��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�K�7�jQѣb��6���>!w���>�_�,���z#O��1���*�������*��l�,��}�V?r4>@G�DM��$��g�T��m���V췧b�yO���B�r��To$�J<�&�h��k}ݟ��ߴ��Sx 'RK�q*:��Q���o�S���H��l���YGBU�3aOM�Ѓ�ܟ��j�m¶�N.������p(Kp+�[���i!4'}�'�8���%���o����0�I6��Jµ`5�h�R��D]�'A�pc���J�sq�`��b���B˽�e�pf��� .�ܻ��a��G�93G	TE�jXȟt-ް;��p�jҐߠ�
��A�5�t̉���G�����3nT�:���P�ټ��|.S��oU�IV�
~i��vT`ELE|2X����=hJgr�R��_:e��g3YÔ��t����% �am��s涭�%@�;M�4�kB�Ico���Id_>��u8}U�&��3m��eQvs�j	|jIW��rE*�3t�࠵�?�%$�;&i��@�@��)����%���'g=!6i4[����
�~f.�I�ⱎd������
S���8Lr��4����lk�#b;"�N�Pĩ�Y�Q� $C�h���{^c��5:9M\�&B��}��d��G��®�5�|^�Ѕ�7��Yͳ�/��+�}�g�"�A��5x�o�n��zY�w���M��������u�t��?�Chc B��ݐ�V�6�$ǟ�v��RC��_� *��w�<�� �dc,�z�U����Q�9��=�G\ŕ���k�z�m��w[/jS�%�fG/�`$g'f�NyO,th�)�MJ��5�M|cw�$�ض�D�:3��1�`p��H�N�τ����-�~��b橀��e;�jq`�����4�������o^b�y�����ߔ/4d��Ӡ"���ߵ���Q���ǁ�ƌ��4��\nVZ5KK�j��������(p�0��7�B@���']�'����w�ڣ�S��j'�(���S��HD���Yt�U�y��L�4�0�K�E���P1�.���DS\RƧ� �(�^�b������A�
�N~���[x�ے��z�#9������6��4��KtO���Wп:�>F�7��ِ����ضl��8U)c
؄ߌ�Kug��*�EMl�R��j>� `�T�1����[`�Q�0��騭�T9̰�
��c�6=�B�ㄲ6<R��n�P�H���bm�`E#�mp'��?��Lg�*��yeŅ��yY+'��,xi��ɒb2�?.���Pa��"����:�=��Zct������ڈ��n�]6�e�n����rN~Y��ޥ8����Ɲ�QA&~�>�-�~��&Ąh��xВ������$^l��N�y�
���[�I�}+y?Y��zU��b�lNr���"��������><���&�� bA��'�)w�����-�S�4� B��<�����jM%��o���y=�^X�A�JoY�S�]�5�������c�62i�ͷf7�f�*8jPj���*�v��c���d$�&�I �~n�}�'�"V���^���2�9ϓp eVX`1E��ovū��M�P�zpX;��v�A"��������q�5"wȟz���\l��-��N9�yV'�
磷�Ӓo����c��'�u�,yj�����h+5�+�N�d��O�ᤘfZ���X��3u����Y=~p��[X����'�T�l��5E���_��-.6ޫ�N�E~ģ0���eW�.����O�4^}~�s��Ez�S�zc��ο�ы�B�P �kgԤF{7^j�|G����'Ld2:��+�g$�
l��z�8Z����f���w VKS��>�a�6��y[�a�dU��0�� ���ؐ�/�S�(��^]	ӳ��ېr���� K�`⧺0C��$G�t�xBl�Oߓ�m��L{*��o�	T�A8�7QI�����"=��A��͵$��`��8�w�2�@�T�Y0�9��f�i������h�v
�$?i��h�yM2_��g�P&
ܚ�ks"BJ�m#F}� K����k{�R�:�T����P/0iZiS	�aT���5��F�ߚ��K��c�)����C8���j+�T�Jp�K��{3~�ϯ���s���M}����1|��LZ�����݀���|��FI����]���ıӶ�᎒9�EF;Blh<�b��5�#�Y(_]A�S@��qx�d6�A��(���%	�c�����77�O8DH�)����������+�6>�Շd&���)f��:���H�C$t_@�St<T��F�dT���&7�k�M������ډ�W��u{���nD�����@�Ke=�]>:���Z�H��0�M~�7��UP�Z����1�0���u�g�mqF�!^���	|V�4"�����_."n�u�z�{V�QRE��z�Q���_�g�C�V��{�y?ׯ����������$�$d)�+}6�[�V>���W��5����E�FWq�3���B+F�2���ޥ�ђ��.�5�T#`*�u]=$y��ۈP�N�(d�R#��q�}�m._B������Jc5�ҳbk��z�N@'f}���}%{�_�ѳ*A[!�L�"��3|FV�)'�)�}V�CZ�_��t�C�V�F��;� �pj2�$�8�<��\��|�j��6=z�".��#k&�	RY�A��[j�`*<�]�"�$Zb��ng��X��]�]V�?�߶VcYpCe� ��d�,���_�Aߊ�v'�L�a9�X��0����!�?kŨ��8|�����p����%���Ξ��y��,�);;^�G��	��Lzx��$�̋�s,|�8�!@�=e�A�JN��g֍��͏����Z��}�Y�)��?@�!y^y���5¨6�5�I��E�6����s�?�.�k��3���"�Ę�sF��t�E��xF"R�����Z����o�1P�}��x�2���E8���C��X�F0K��8+���t�\��)?X�v��)�WA�UO�U�(&3���i��f���K?Y-ڎ��;�a�?	k�7�I&I��3\w������
B�������5<��wF���iDF��]"t���&j�����z,��
�S'96߇[�(	ԗJ����T�Z���*���CF�|%0��;~B���2���*[ѤC��*�{����O_��V;e����[r���	Ӌ�s���g����ao�T }f��-�91/�{J$����ñ���w.�!�M*h�5�<�	:i'd"��X�;4a���b�s�5�&!�0��|>Y&��e� LŨ�4I�R������(�d%�h��u�91�5��R ��6���p���M�z����p�'�����?`�Q6C�ʛ��m�V���Z�	�������e���C�y�� ?������|��b���|��w�&h�d�aA��/��EU�8����ѐJ��`��0��������T #�-�]L8>�9�&_��T����2D���U�ܛ����p��׽o:}�iCu���Ή���+v��R����&�\�#�Jv�x�,x�5a�:g�W� j���	2yq�;��'������=��R!����2���	a�O�L$���Q��#�W�
#�7��B]�/d��wt>�}P~*$�����7�5LT��N�~��\�qF]��#�j��p��� ��B��ҭXѝ��p�K�)�����P�Z	��	��Z�)�R���vR{�3*��;�m+�o�\[Qx�j�.�bN�:��.OB,������ 3Z'͌�&�
���NJ��+��o)T�,��4���U��A���T�r�4`����_H|�#	��佹��?߬��-6'�7�spZ4=�N��9�J~
�'"��]�]���Z%��a/*0�mv�X�v,h����P 
b����T.� 's�gJ�Ef�(MLN�S��lW�5�	���O*�('܇g=�*G�+��ڌ��Y+6���\�#E_�CWY��T���T;_���;6�6��>�=+4h���w�>,�IÔ<�'�u�+�#4���_�%��[^��롰2��J�݌��w��آ�N��\�R�I��ͼ�E�	Ҽ���n��ُ+�?�T����j�<,��w�(���3`���W��ҦN��M]Ig �����n��d`D��6�����I��d���]����A2v��`/�rZ[��P�;�]fD��%�?��2J�2�nҢ���:�c��RDDg������}>�L��dO�L�褤[dgd5%C.��z/�7i��Vߚ+�{)6��	��V����8EK�>�?�?b2�pge�����FGUg�nK�w4"_�����P)�nͲ�ha�`3t�&%���M#����1:d�z��'�����q����P�Q̆��u�bU�"��-<�֏��	����زs��a#�ԓ�q^��`�Xƭ?�+�..���`h8|�|��Q�bJ��Fj;c|���i^��/���C��G��6w��a���#��\Ԑ�x�S�;�|������*�>	��沈���|��8�q
����X�R��N\=lGm$�U�k�(�"�pصK;И�6�SB�, _b3�ƽwϛ�=-���g�ᱥ-�]�x�����(�Ŝ]�7�T#�L@1����@����I����!X(�5d
C(�����sV��tU �<�b(\�І�� }�\��[ɯۈJ�H|=c`�,N�Rk��9� ���-u�8��jB�;��[��ٍ�%�Φ=U{)���#U(��"9��ӷ��9o!���8�ϒ
b����9͑���vag��z^1�T	�ͳi��Y�ni�o5����⻅�Ȑ{��x��4A6��< �h�h�0�,��jd���Q/I�̏E��WP��$�?�ak�=�[���!���5���"�^��m����јʛ�ļGy�5�)?��3�K���l�)>AEb��R��+����w6��%�a���E�Bo y����0�fi�	�$@��}�UgV9q����s�)�ƥ�֨�on� �˒~��Rݳ���ݖ��`Xf@�_�M�ڣ��ʼ���T��Ֆt@�/h��4Xw^��q��#<3�$)��\��j
*����xֿ 4ȾL""9+ՙ���a�.@�x�&���b�����,?����;DŨ�>-�요;��\�l"�l�)��M
�k�f�-���J*�N/����m��Վ�㹚L�+W=C5֤M�:on�o5zw�����Z��\���nl�z>��	0KO	zMH� >�8]�Q�/�?�����(t5<�LZ��Ey�w���G߿l�bԂ*�3��]��:��ɒ��=  Uom�58�e;�u���΀�i��/�D���$@cs{k�����?ݛ�euȘ��f��=O�-�k���h�?�Ar�����N���
�_�zNά��(�D������́8�>7S�����QR\�M:�uʅ��C�n�s�Mį�sR0�����%��Q��u�2'{�^�b$��>�t�jIm�7���d��l��>���^z��x����6��}�O2���,ת88�J��e�U;�y�dL81Q�z�c$薱���"��);DN��Y��ߧY�n%ȷ�3Qp��^�.����JA26dC�����"n�6���U�1s|���S��i&�r��LU��;>��0�̞!5 �O����vau��xh�&Ү:�j2G':�u���a����������I��=��	�XAh��f�:X�G\�@y"ž�aNe�s�(!I��z�U�s=�hȭ#;}s�����j�?��_��u۔�-1n���yAk�Q;ZZ�#BHъ�l	����T�&w���6��k�:� �����v�Ɏx�|eP!d\�<๳\1��e�5Cp�WI�I�K�C=����4/�� ���� m8	k���2�|+���r���G�"DL��+�V�y-j��|��0&Q��2%G�`!����}�N ��Bz`ޥ����ڡ�Cr�]� �� ��{��ͭbA�9�z�  �]D�Z�nc�aL_e���]�~'6�~��us[H�����g
��S�φ� u�M���f�#��h*����g��.���k��o5Wn�Q�he�;�}�w��L��`�ҵ�EѮ��Ғ͑��� �ށ.rb���j�~>��eD�.�T+�0u	���o��c����`����������1�$'��н/]��wi$i� GNg�?�,v�<C�me���1)�}j\�N ���m6�;�9v˥�ZY��_�h��ȍk����w: ����СOn���-S9/����|r��ov��}yuWf�F��y%Q ��Þ���蘙A*���	Qb���~��8KJ��݈bO��a*�4�� AL���;%/K��[b��"����q����:Bh��p�2���� �a��&$���28 @|~��Q��]?H� �,h�lm�9��W6�Ym0H�2�5Fi|bE;��Gv�).?)�@K�O����O��zH�`�T���R1s;R�]YW9�jI��/=6���Z����Y�F���F�rv�K�8�$���U�������Q��IrhF�������tQ�'���:�B/�|d�Ax�s�
�5�Ʈ�}fB-�E7h��Ė��T�����y-޴d��%�52���p߮���Mch�͋�χ5hm%�޸��6�J����
�&�*:�e�W�	�������Aӻ�B��b�aǺX51+�d�����ĥ��"�(m��)6K��6�f��O�@��S�i�ڥ���v)l�q�P(��ݒ~�F����b��Zl�ex��'���.3%N{�ᠪK�Ŭ���_ļX�93.cz��T�J��?)�~���������=30�x�Si������ȍ����R�PO��C���׋�6�0�0:�徃*��牤��r��l/�55ύ����Ǚl���
�=�xǭ̽GH�8�?[�1x>y�2�8����V-� �}��iB�f�1//�!�dQ7�?,�WWP@��(�S !���h����{<	Lގ��-����u̅/\�!�:��_�}�O���?�>�F��ꥀM�.��?��������t �y�?���#�eϤ1�؈%ʬ�L�ݗ�cM��]���x�c*)��U�g��O�5uD�o��R�uk6� +y2�,�	�~>>�Ϩv������>�z���e��'�w�K�c	%J�'?	P��
�>#�]q���si�d���M���h�6X���?���qZ��!���X�q=\���0�)3��ɍn��3�+3
����l�_�I�ee�ꌥ}�0��n�1@�0�z�]?�AS�˼GVK�պ'W,��eaha�VΙ�������r���n�E��`�	զ�//��:���&󕡯��w��(��z!�Ƃ·}�A]����m$��NZ���M7#�)��dR�(������+����t�i0�P�ɟ|��M1���>�7�}{ 0�}I�����?���ț�ABG��6�S�Q���������/�f
���W�8�q��`�'{��]��y����ί�B�"�\2�F��g��m&p̕#�}(uc�~
(�����$W�ќo39��lV��`��D���Α\ԯ�-���4<=�i ������Jv_؟R��@��=�=H�V�`��5[t���i�"�{���`zKh���-�'�5�:%��v�ݠ���hL�k���S�3�F1�xswL��8���dB���&$��Z����Q4�$<Z>��m���w�H��8�s����Ȃ��������&�GeÁ�� .)Sw�ͮuC�
�p�G���!�!|�p��>��r^�XL;�j3o�-�IV52�O&}Y�`m���$�o�	SD���\�Af�>�5!VF�4]|<m�gC<�AR�"V (b4Y�$��}��J�7�ݕ��o�[�9_��y��w��~��&.]�a���_�iUX똴��M�C�����1��g'|өJ��8?�Z>4ӯ�v��V���)f�<���f&���|����݌}Bz;�#l��Ҝ��A`��O�Z��MY�����@צxǜ�NA�n�<gU����j�c�#|!��(�c�
t|���$9+U�
�Z��ɝ}�r$1=R�*g���������֧�kQ�Υ�(�����[�����q1�s�e��c��W����PÕ�ً��5��Y�mP 7_wX���R@��5 W�͋ ���>3?��1Ar��<�QL�2�;�h(Z ���s$�e�"���=�B��8^E�/�-��ZRᠻ+ B��i��8�?��J�o�%=�Yl��@�1��(:=�wDh�R�4�_�aK�$�߯�dM�|���k�
�Wƶ�۳)Ӝ�P{�c֌k��m	����+��~PtK����&<��4�6��f�x�������9��O}iS"�#h����S3�(��	b��� ���ԏ��&�#3V�QK��o��'p�&�T��㤏[v��� �-�7�J��9O�t.§���19�Өǭ�^���B!��y���J9O+��4��Ò.�%o��Y��`T�2RMP_�7)�k��ZR�jg������S�W�u��G(������s��*��-Ik�Pο�|��ٜ������͌���r�K_P�|��ԫt���w��iF�`�NF�����)���4Q.}��~D���"��u�g&���n��qx`��q�����g\kj'F�DGX`�D�P�R��Z�|����H�S�H��<�u|�U���ЛN��?ѣ:_�V�4�[�g�t*��w���VN,i��~2%�Y��a�B_�,ϒ�V"�/!ihR�m�%���M�pA����Jh������q!^��y&P'�7%TM��Dm�b�v�?�{8꧃�GJr(����+���h���LH�\20�ĊE|�S���r]����Ϻ
"�����.��Vi�tJ����zK����-���%�F+Lc�5��t���s���+��w%���*)W�LYh�R��M���T�����m+Mn��,�R�����(�Rʹ��c4�ڂ���̻XN�����TQ�A�b�#D�L��ހ���Э������J6fXjK�A@d�)�w����2i�4�����A�kJ�b���]���|}�����ꭾCK/����O�,_F�I�\-i.?c����J�&�]����2�w�"���|���Y�P�T�N����X�ع��%u��s]��N�Q⾗!+���^Dh,[�tØR�~�ٞ�K;��w�J[s.ڷ���
>X=Q�D
�g�[`�y�3'�A���"]Y��j۷8�Ǝ2������|:%i���#�EY��qY[����T�&�X�f�M�?ʡ�bݳҝ3�%_�FД��0L��_�}ڋ�ۅ��W�\��di�{�TC!Da�n���M��R[��z�P2�* e�������*u�����	4��G
���-TOp�Pv����@�x]��Z�5Q��̿�pLgz�E�>�Q)�	.�1�'M�������j^��Mm�d��ںSZ���\LQ���ͨ������y_��=��D�g	$B-Rm|/��l����f�vOi���z���	^�2�o�����
iT���{�:l����_�ֳ��D� {��X"K�3WE:o4��`թ�)�5\�x��B�B,XE�RJ�L\���g�I~�&T~���IU��QNBW�#���y�y2LH�W��������ޙ��x�f��Y�"s2�Ry�2�&�q�I����ͨ���q�H6xm$�:n1�$!p��I z�t��W %�eR��@���d����+��u���P�S�1�pV{8f(.ܶk�t���� �5��Y����z�*������n|���J�Nы�}�-��u>�Q��pZW�ؐ䲺�G��hL�4��;2Kn2wYOvga���pl��r���ϱ �J)��~��>M����X��t�V��D�pe(-M�ӱ��-��w�)9�<g2�qmψ9;��ʳn���f�&Q�#01t3 �����q~��,z�����N�
D�D�,����O���.��/Z%BF���=:�f��u�2���"��̿����M�k\rT�l9+ra����Z���.���"��}��d���k����4�W��������Eсfj�*�$�Ի��k�r+���|��dig��g�/}"ؗ~�ۣ�Ztt��+0��}(Vm�C�E��hd�>��PG���h�g� ��9t�x�t+�}r��3G���%l� q-��ޥ]�s_��>��L���n��ۗ�A�9P����k�푩� E�#�L�w\N�g޼'1������ښ��^�@
Ú�-메_6���av��Y0[Pc�
��۰ヂ�� ������9EY?"	*��<�*�Q�!�CO�O��+"gEZ��{~���3-��D�yMcd�O{	} �͂$�M�/��k��߰�=d��^�m�1"��@0Y������.$r�� �R���=�*�rw6�(}�YX
l��eC�m�)����G��G����g�QNv�е#�<9,|�:F?�-���΢b����TƲ;��p_�|�Q�J�.K�<^_}q!�L�x��ur-��w����fo�#��nS���=���H��,!�P<l�_h �067l�p���z�K� 0n�Q1����|e�SC�cD�ϱ�u�ݱ�f|�Gy��.�Ea�U��v�N�B���,��۳j�k�p��z�a���jR��fx|��1;*�a����m��RR[�pB���d��}��a�T}���>OV�\�[�[��0#����y��H�1mի,d�*8�K�Qϐ��i�s�%L^uY�z�>%'xX�sG"\l�R�CÏE�fՇ�	�-ҙNUi��������@�m~�P�ǞX{���	%GΦy;%hK��zUC6m���jh��
Kπ�e���.��hwBm�}b��`�*�hޗ�S��
����Wb ��v�E���9nB=~ߠ���C��y0�@���N"�N+��kT�E����t��;���6���<�:n�mYõN���`�i��das]V�&��3�'{:���lG�27e-�H��E�l^����W�TR����w�Q�mI�`��#\OL'�/�͌��Y�Ɯ�}�UE�b�B8�ށ�/h5薕�{����O2��� }J5�9Qnu#�����D{���-����'����Ḇ�7s�qI� 9Mn���:5�͑�`I4-z_Xr�=|�p����#\iq0TR�4�?\H�:���ς�n'.�N�{ji��%���=9=��	M��d�!�-M��ӑ�-#'2&��Z�A�IY%AT�!���`��^��a� �{dM�]�J�����V�_AO���A#��e'7T��f��%�.�-*���c��W2��躆t���Awp9���f�J�k�|�W2F�5��M��*ke޺�*�+�A ���7��\���c�
�.�������B4��
��zF&ȕa�^����N���:S�B`X]�4�`~���N�cS�f茟68p&����j��G�>� !���w�M��#�I���I�Z��E�/m�y�����W��pχƈ�8�z��UM�oVF��{��)�%�*�"������������.�Y��=�{�tM��.�z�[F� 8�AomrH��$7�j8�=C3;U,��Vq�a9�����M��<���T�� k<�T�0��\�zo'9���	=���JJzj��:90J��[H_�،)�>�{q.��~�g!�r�r��KRO%���){:V15UܮZ��w�7��k�9�o� Y���BN��87 )��܀C��A|[�߽^�+�A���$���8u����j��7���ϴ�Jh-X����ɸ�C7�^< _~��|e{�W���]�7I>ԝ�M� �PZ�tB�`$�iN96:`���
&A�px~�D�m�T^l`_E����FW49�6t�A�4<���ǥ��é~�F0̿ѝ���
�.b���<�[��jR�p'%$�B�!v�Y|��@��b���r�Z|V��P-��%���^&=�s��F�9%70)��L,��O/��r������Sv1}& ��_��Z4�-�*E��gT���k���WO�=9jn����|�XZ���zn�U%�L����f�;F4�<�3��C���g�4���erl|���x���DUц3Y�'��c������h��Hw��|��a�O�]���
�,����wҡL����l7������_{�ߴzP��$��^�T1�i�G�Q��Ѻ	���f� |��2?��}l��c�*3#7^P���V{���\qm'uRg;��ЪEﾜ��b���}A4_y`����T��r)<K��q H� ��ǰ.ݡ0B�c��&�������ކs��祤�mMU;�s�����	,��B������p7{� H=�L�v���k����qȓFx�)B�E�OH���L��ť*(xD�ű�-����M���U1J-��`���164ƫd�NQ���-P��m�ȉ`:s�9L�2�d-�H�v�;�;�V�e"�	��c�s��L�&T������Q;�`�9���]=LS�x-�1G)ʴ����r~�B����u�1������O�)n�]���b��G֭?���cȨ���\��k�Z�giY>�#�={��v�h�n^�����.UTL %�RU��k�dLɥe�^�VWS���_|�͈���',d�>���>���Nߪᙔ+�P͈�jȭSD&�X_�寽���%�?�V����f>ץ�EΗ/
��gNٯ�����R:�jJQۻQ�O��$�`�^5�R��")
�$�n�͊��?�ٮ�siP���7��/e&����ֻ����>�/}x��E�b���vwb���i�ubM$��U7�)��ald�n�
�2NR�F�܃?xWm��|o	9��cO{��D��9�j��-\��!G�v_��*�Aަ�߾E8գ�|3c���;VJ E��q��v�y"�,OS�}��i�L��I����TL���ɯ��(|�n��I���U�I���{��(	��Y�gL��������R�_��F��[Ӑ���|g�%m-��SJ3~�İ�Y݉
Eψϭ�p��eR��k.ɠ���g�`pJHm$�����Q1:��Q��Q�9��Ss�LI�M��[�)S�@��) ��̱)m��DL6DDs9�z��N��M�$��mX5�
���oM��p���	EYa�����3� ��qӹO����|e_
Sb��,�����E��ry��59�g�3=�I�c��)Et�[�)c���sh�-����ޒ�toa�bd�0��GSzְ7N�M$R�|�����͡��")*�t�|�d�tӁ<�����z�b�����9n\�k���!3g֫�@$��tB���M͌��B��=<��� �5F��i0]D<�ް[(1�$(Ѓ.�S�L�5��l�j����1p����Q�V��s뿓s=xt5�.�̘[��b!�%>K5��Z���.g!��3�_��d}���8�jH_4"g��<w�ԗ��xv�J���"�!a��;BS�;��������Y����@�F���=H�Fh�B' ZMkcpE���C�z��:$8Lc$g����;���Tbh�ެ��K:����?�#nI�D� Eʐ	�n邡4���hy�X�c�����U�
���:K��7�˹?JǞ(�5�/ ����ҏ�,Gf(���$�*��m�"������K \⃳3�3�;?S��!��>��U�M�,��ا�v��؟��yK�e��$+����L�u�{G��c3���"�$3k�l��+�H��<R�
����3X_x:{8�Ėx���	��씲�yu��^=�2��L���?�X�d�͛�z=|�Dr�B����|dB�lb 褲�h�N�����G�ywX�E��� �h4���QVX0.:��W�T���<j:��k�^�b��4�C�Ò}lrev�7�M�?g����)y���d���e��1<�Xb?3�( �G�]��H�\w�=�����yi�SX��b|i�q�t�����y��ˣ:QE⎺_	����0If@����W˺��
�����x�_И~zƟ����~#q�>����T�W�Ls�E�n@.^O��Jp]���Dn��p&��%�7��V՜�s��{��3��3Y.n���2�VWL˺�NWt؄�� q�xr�갩���d$���c��s� u�I���;$6���j�<�c"�^N��������i�E�4Z��M��Q����/�W�mU�MOu�<d���7%��vq$~Լ��J���q�� [�#4��*�n���"��|��V�)���&��*��ퟩ庤 ��m+���@�Y-�e�
a�@�J� ݿ�_B��<!�+N��ld��Oa���뿩L���S�4���uT\���������ڢ��a�!����%Ƙ��	R!����<$���#���JZJ,w'I	�G�8y"�-���~�gsu=�櫙�%c,i�y����Y�ոvGZ�� U��1|��	��@g��S�3��T8-�7��-��`�c��6�^g�f�DCR͌�/?��;������]/+����B�K�Sre(H|�A3�������{��$	�v�p#�Ǿ��ve8i�yeOs��P����s�5;.�o$��6{�IzY�=�)��L�G�~��Z��C�G���]�Q� ���|8��OpQ}�j��m3�u�����(W�D��0f�x��".������ɰ!�H;�H*�_%h#��l=�4S�u��&ѿ�2ю)��Կ������3mO�h*E�l��*.��V�HR;�d�2� �R��e����'dOj���@��7C��RA�i��Yc}�Dc/�a��(q.��c=�� 0��Jl�7ui�Ϟ'��,��R�b)T0��E�7��^+82�N�Rj�#�wm��	8<3�7Z��2���x�ڋ�tT����k�ȳ�oY8PJͰ|9U�@m�\�����p0\d�6���+��k	�JW�vP��i��o��#� 4�ԗq�KO��L�6`�q�52�������m��m��-nü�j�W�&+�˚�+�M�����OU�ଇ(��5�c�:HZvXZ#E�z�ʱ:����T-��7΢���� b�@j��7�p�<��7� ��MP^�y�J��z�]p���&��S����<B��|�G����s�Z��qN��X��R�5����]~��Ǐ\2+%!�+	�q�paf�k[�1|�0+���8T�;��U����x���EmA�FG�v$c/w���NtNq��v��1���"ΰ0If{͵�	�х*���y�ZԵ޵HR2>D�-x�k��F5,?m��aX���x��9c��b,�1�R���2��kr{FR��;����iV��սV�DD�Ti������3����K�NC?�b�\l�mDRd�)�M��ve�y�@H�\����Y��OO~��ւ�!�� V����EKA����n�wIwS�x3��?��_�^0���]�n�7n���;7k+��}�5'TRʆ8՟樇bN�#�T_�p�gǩF�>gP5�iMR����?3�fN�m��Z��`'.�㼭�g��az��HP�,t��X�GB���Y�%E���WD�hwx6�N
+�~4~��Z�7kv�N_�t1�g�
�@8J��v��ݮX#�PgS�7T�A㋨A�"}�$NL����}4�&̄�q��M�(?V�
{�8-'ʛ�e<A�{�IPn� H1xk���=�w�
�����?��G��M-t8�k�R��>��ņQ�C�h�K��N��M'e�l��  h�K!�\�G�=~l��x���۴5:)p��6�y���(�0���w~��u5��z�D4_|Y��%�?!$�]e:�z�Ez�������bL�|���KHrw�
�C�"�{�'��_�P�zTA��EBA��z�%�稉MD��v���j���oXI ~�dP']0��g�����
��V���IOW��G-Dn�����?��ÔW�;T���k�� �1Y�o7�x��D "o,tK��]
�mw�������(�U�m�oky�����R��������� �����eL�c �|��A����Nr%�-v�לH�I�o��̋���.���]�Ҝ��,f������'��M�����^|X'��n1����7���XP��@+¸��D>)�2x!.?3;ep�.N�d�~X��ٛ޾�&5��V�!?e2!�M�I�dS��&{�
����G �����l�+]��6��:m����Dv�|_m�L��kV�,�N�%��G��kl�T�۸\g�@s@��L��)y�/�X����6Zc��kt��1��|LR�0L9�`#�oD�os����@��KT�ѭx��Q���hV�?ѷ8�z�����mG��b��*y�+t�5���>�eE�M	���v�v}������Q�,��Q���5�5��`��OQ�4cB���(X�����C�oNY��i]�������� ��g��{��Q��h���r2�k�Ahl�:Ux~�B!�)���6r)����Mp&epJM��	S����?Y��Y�����Z@f�A/0���)��!L���-�#k~+�Yc���2̅�7~.;�����R��g���.m���R�Z��$��N\hY�qVK�g���zSe�qV���ҟe��E}6I�[��O;�Н
��.K�~|ۈ��`4�+���E�,c���`D�y\5���fSߘ^sy�)8�RFVϭ��+�A�m�����fö�k��
����}g'˸�Z����	uה������lZ4❇�_�8z�
�tH��.���.ۚnCz��0�=a-�����	ː�B:^K��t���=K#9�@âA�ѡ���Q��br�`�a^����<`��Jig�h���xzz÷�c����[P����wkGo1��g�hL=�� �7YL�0��#�3{u�3x����&���\	j0,��j_ %Np!d�w�G�i�N�#��� ��&��2#�X�yUQ�C:���[7_n�3 =�A�Hv���@f��U������au�,<R0$!;�`�\o)���&���|�2�P���KO,U��>�5;�#J�r�2�_�Jw�]�}�f�z��p&�:rQ�ܿ:z�(Us�������1�� ��Z_��f��%$��NN}`L�0��{v�i�t?�{`n+�2J6[g2:�:F3���.���k�h6���M=h)�@��s���S�h.8�Y;0&�ST�h��ZΉ���Nk��K�� ��v�$�o6�� � ��.�����֬�/��Ժ����s��i��M)~t?�/��	����O��� �V0
Z��e����y�w��l�� �s�y��|j�a�����"s2� I~��S���}�*��X5�AZ�Y�@sX��_�mnO�R��\��-G�?*��hyL�}�OdXKm�>4��i�("��Fl�A-�&�7��μ�F{� g���M:�<��VҌs[T�\��}i����`c��:���~�Y����2>qH�ͯ��7��X���� (��>X�>��j:�@fd��kiY��wb]'�Q��pRc� >:�Q�����5�PˌqP/4i^���P�]�;����"օ|�r��c�T� ��y.���/������=�K����y³�-�n�[D���칼�
�~J
��jj��|�j4�xk'��U&�p�A7����B t��у*��G@�!���O!��w��A��
��ˎo�Oxi���UüI2B~;H_ְ(&�dK���ً!-W�G��`��@��5�Zc�O'x���]�8�@tsV�ݫ>�n�w����N��.:�*������v��]h@�Lz#B�]�Kع#��D���*�9��TM�w����IM͖L2,��
����Ζt��w�$����M��&Q	��a�FF�ȥ	��b�Q����D=�f��E+ޚ�$�������P�"�13=Qܬ���?>���%`���?�}�=CJ�٥p�C?vZE0&��7��1.�3$U<�[�"�>[���4#�nB����e��P�w�����&|�b
xR�bQ.�ڶaS$��u�����$W(�cCn�k��%�-e�2x��$L��Y�:����{��y)qLژ�l<V\h�;���K82ߕ%�#�|8��ԤO%�m�躪.�=�sF����d�=�6��sҷ|cc�,ǒ�Ŋ|�%iX�<���#F&w�zQ���o�nye[�a��H �*h�yS�Ci$ĺZ����f	�\�9�ݵ�$a|��#�k��b2 7QM���]�ƥ�W�T�!0�5h}���:��\a�E�BwF��0��<�ۗ��ʉz���"�S�s��o@[����	�A3I@tS�tQ��J�MC���f��+9���57�m��?Kav�x��g��o?�յI�~9u��0 R��'�=ȫ7>fc�g�ə����)���w1qi���n{A�p_��P�F��M��<h�i�Ӧ¨�Oʰ��]�3|,�s�3������9�n����-���n���OF;��e�C�}�Mi#x��ȪBV��2�I��I�����=�;|���o����.���*�`�&����341L��n���ZR��ͧ��#
���d+��X0
ԟ�6��M�<�f4��ַf�y3w�yμ~N�t�� w�(V:{/xݺ���C�R�4��εFE,�#]�&��d��`�r��̆�Z?7�Vy.}������g� ��:W~Y#�O�S���:$%��4(y�<���ShY���t�P V�$Fm��q5xcM��V�g���wOр�K��~���j���@����T�`�Jn��^v�3n7�B�-�E��a�	jf���R$V���3j��<���͕`f&DY��;h;��tj���H�q	BF���? ��b�{�>=p��X�!�K��-�2W4#d��
�^*�;��k?	ѯ�f���͏�t��I���.�5�X���B�Y�l�=V���8K	c��39_�JH�ƼsBn�ě�W�K1�L	�t>�FY� B�w�����5���'�5���}!�pb\wy�z�Y2����G��B[����ԅU�F|���)rP[���"S�Yݡ_���.l��]�1ruC8�=�3�և'k�F~�	��+���yNdylPcR*y��l�l�� #�l��a."�w^R�ھ�����u����92s�����9��NfF�(�x��a�:Q�!�J��� �q�t@�E1��1~ںz�K�/,���]��HL
Z�����YW��O����9�}:�m��bȊ[,\�R�M^�o�*���p��P$�����"vu��{���2�\��8>��4fEr�8�.@g$��6ω�}v7�7`i{+g��'��E�;�1��2���ܿ:\���e=��M1�v�CS��Ӫ!p/�<�p���-��ځ.�ux�l�1j4�sVT��֭O�0���s��\�PP pI��j@J�z�����3v�}Ě�'�Hҍ���?�g�pWII�0�a0���h�{��7����r�Ԫe�@�[�l6?�o�	�h�#~IU5\
�g	$�}C���j=� ��!�ۤ��+��ޓ�榃�rƥe$A�L�u���H̙1���$4��F"J�ᝬ�C�gGR[(��C�Z8mJE��Kw�L�u�f�%�C�w%��\1���1�W�n��-�.,�GJ��	B�hj�Q��-�U�"���S\���W�Tr��[N"P8>	PY�#'�Y��L�W�d��d8������=c�z?�_� �=�
]�TTeНBaا��I�>��#����418Bn������x�����w�_���Ӑ��'�j0)U/�t�&��ݕB����/8��o���lج8rFEa�1���c������8�Y%�bͨ���Հ��-����G��r�`C,��;<K.!,6. ��N��$�`�C3ß1� _��S�gF�md&�>��Ρ8K��{�S��Ԕ ��Ҧ���vJ��3���	�V�Ԭ��ev�28�2�G��;�����k��I�8�hEC�ȥ��H�����1 �6O�������_3�GYF�QBz*�~�BNh����8�-F��",�W����b��P4Ls�i�Ƃ�a�C�_���	�ƞ�=���:\��*��c
��Q�]=S��r;�����z������Df뫣s0�/b���pN�Q��x��b/�|ֳu���$�w�`���k,:}9%d^(�KVჾ�X��p:��0�1��r����׶�^;����8��x��:
A�hK���ճ��nS~��>9;_�D�6I�\���V��C��D�R�M*nL E'�{␡��/{L3p-���9BQ2�,���o�����+&|�Jɂw:����V]������0��*�����m��P�w�?=Qۗ)��X�����&ܞ-�)YPK5Y5/]���㶡'z�>fN���e�������k8W(�x�97���:S��;nj5_�M\�������Z5��Yn�.�!J�/��&*���f��~�G4�Ղ�������y%�����5�b������<訙}	u}��>�ͦC��K�k�+�#�G<�m�XL���:ed�2��0��lT�&�ҙ�b�7�]�qJ��ڣA�j��9>ρnsL 
T�hBM��!z���$]\���;?�0kIK�KQn���� XR@�� Z�f�"�Cf7�X迺�F�S�bB�1ri��R���nj�\2������͒�ȺQ;YvUf*�'L{�c؛}.0�g�9�
��Q#�0��%�xH^u�My��y�9ܭ�H�v@o����G�xLh	#כPͳ��m�"�� K�9�p�)8*-����n�2	c�`�yl�N����S�N
� ��{�Æ\
��*��93eIjs5�]�P:U��H[35vu�r�Z�X��zE�h]��e"!�R�~�s	�ȇ̦Z�7��"��Ո��\7�@���D*c8.3uWQm���^�;K������=�6t�\���~"xyUf�~�I`���`O� �f iy�*�s�~���-.��$����gV��/\L?]x#f�ҳ�[tL�ٓ�};*x�P��K�e
��_�mh�)��0Cɦ<3D�;�opU�.���z��Lm����7	q�}��(��A/t�.dh~�m���}�D��-�O��������O&���*�~j�[8�#����G��[��5�����>���H���(SJ���5�z��.���bMOe��>p��"�D���ʂ���]6w�W�Ʀ�Sɛ�]~����Q�r��&$��;�BRI����&�/����-�pϢFꇵ�	�S��Z��M;���s�s+�9.�X��K�����}�s���[�dZ5r�|ġt�C$qR��}:�4hR��YNlL%��	z�1�;o��K/�����N3�����^�xn�k�w�Yx�lCܜ�M��b��2D��z�b��U��d��QÆ\F&��p���S�i����A�����gM��
�6B�� j�ِ��U8��c���:=lԭ�J�nH��aӸD<�k�tf��R�bG�;Y(x�)�Db
/�L�K_z��e��������͂h�r�Q�`�:j\���\�6.�1�N)sp��Bz-�-|/�6�ҙ��\��}�Lo@�I@	x�Y��i;G��G5�K��������tO�9�%<dCv�ZCs�X�u>!<z�IH<��#�t��UZ\��B1�XD���#~�޼��M(�;��J����	A�|�N(k�-�Lzҩ�;c�X��鎏4��*��mg��<���m�H�P]�i�����+��&�����4%C$=b��<��� w i�'�8~M`X}�[q�����	}���v�j��w�[�*abHe�CɆ� R' �$�xkj3���Eu39�3,l����,[��$�Ɗ�wv�;�L� ���!�.�@�	W�]��~�<8�� ���-r p9yfU!t����"ו��,���O�t�> =�8�I��2de�a�V��� ���N�e���a�2���.�IJ���e��]�Q�8U�"�1�D�h�_��F��h¡!�/F��|<�TBkdL.�y����Q�)��a�2/�MsUb��x��.�0`x�T�>r�6��2@u�q�Ԅ�=~i&�Ѕ�	3 �)9V9�i���»%p�Ǔo?�I�E<��S�ٴ<���h�h��f��8a��p�0!�©���ΠWI�x��l*�rR�AY��, 1�`P]�##T�JB�x�x!͠pl$��<IO˒����a,�����솉���$Xo��߰�r�vi ���!�YA�����.-��q�P�=��^�0��Iyע�1�����mz=����[RJ�������ROK�.�I����N't�n��q�]���(49�U�g���Q=�B��qȳR�+pR�p�<2�is�t��#6�Y[�Z�u�<���{��$^)3��d�qF��D生�PΕ�ZՏ�������k��P>˨ޏ~F��	���:~)�@���Ř������_�,���k>�l���e�VT�Ԉ�X)�J8�b�N����y^%�t�p��J���R�-mU��#l�C��2h6���&C-���J�5V;Zm2ocP���`u<���ڇ)�Z�2��4S�3d<���M7c��[�������J$�5A����*U��C�q�^�	qk�����& ��=�*f��,,�T
��	GΖ����m�J�@�X2|gi��^IUYiM	-O>�|/A��2�TB�+�L���2���(�e�t��9 �_����C=��r"��$?˝׉8��14N�*�d\���+On�=�JV*� j�R�K��s����� �sGY\�s��h�_g�K$Nk����Աɦ�#h!?��J<{K�V�I�&�w��D��Hm�1�� 
���^���<R�	�D��� �ޡ��&>�*�����Py���xCA,��e0��J?�Y)����Q�|(P��-�o��Jd\�,p�-7���1,��l����ԕ��Y�����a;!�5\�q��ӿWZ��q�^]%c�����l���8Lڜ/|����oFc��ܺ8��7Y��q�r�1��)��hB {�3aQg�TR��ދv8�qf��=�6M�LJ.������@р�lu�~
�y_GQ���_
-	2��)�p��&.�륍���ۗs��C���`�<�k��ږ�����ݚ}�&#�>r�cT�@�V����C�dqr{Rd�����̈́G=S��Y{�`F�gp�h���d"-L��x�ѐO��l�%��$�+70���'B4Ռi'&�5Ӿ��uTRl��	x��I��^�Tջ�/k&X�*�*��VׇDNr��6���3r�U�V�>?������x��|�uٝ��� '��~����6�f�dõ�6P)�����6A�q;���B�AX�}ug����e����cS��YP�s���r�H`����A��~�E��~(%L<\Z]������Bv��k`+;ŇeF���V�([��2/�B�#& K{���Ze#?\=S2s�:�c0��"��	��W����*��g���{0���\�&^}�_�&���~L͹1�C5ɞ]�ȇ9c$/�2}9��?�}�0�*^�| �1��4��y��MF�=�9�8N��y����F��bk�&���@���
RBj}%�˱%<使X�	�\��wn+��ƸNK�u�D"��vO2Y��	J>ghA�����>�W�>/t�[�P�8���䜮�n=�qv��
'ud㑺6Al�6I}����	MI*��{����z�=����)O�x���^�����ڡ��wr/�;���ئ�h鮜�m��Heo���l�>�u
�vO�����٦pFq5�o��+��ja�'��R���.�PD���R&�U�����:nN��e��n�I�R���2��^��l�f�NચN9Q�G�d"8���S�(x���ȄO�"�����0�O(4�Wd�
��$Q�q}��R%ny�R�A_�H�Z���5�K	�H��Oaz�XH&�"������J���b��lJ�/D{(��Ț�@�G3�������%Sxz�V��,ب�����L[`�b:N��꒕��",��0���b�����e�u<���
u��=�fy�B��lW��R?@曜��#�ΐ �h��G\�eZEa�ƣC�����}~��, ��Ĵ�HI	H�h��MY�:�ID����
���a_��%W�A~�/�O�}}����b���>RQ|�:��Ȝ K�~�����G*�DM�o�	G�%��Oy�D�8��,��QK�Fdl���4���/���B�������*�����໽��7c���n��#oL�V�ʉ���{�P�QQ��OD�8�!tU��@ �P��ʳt{	���Ũ�c̍���,�kwx��?9yp��=�Na� �Cm�����*,���>�y|\(�%�@7�Q)$<����VHK�ܯ8�apN_`��������c[nPqz~�������L&&EYx�g��wB��4��,�6xU阑l���n�שc�3j�gL
<1��Ka����~5���gI�1��p��]�xr����5��u	��G�C�
���k�aS��c��8�
�*D�zk�Xɠ��r��1_�E��%
��5�Z�s�O�H#�>��� 4z��IL�����d����^�m��R�$�ݕ��	Ų�6��|W�l���=m&bʣ���D�m:��&�7�.�J��B+:ɯQA�f�ȮtU���r�K0-տf�q��=��b@g�g�Z{��i���B������W~��	6־��P��GKo��X�`�-���M��&�����	�;��*jX}5tƾٝ��3�U̹�[{sGATe��;L!�c-2Q�����\������
���j嬅v)������&J�}m�8澥A�	�p��� z������b_�t�")J���KtߥתM�ޝ�?B����I�Ђ�:6:���Z��:�W�F��7�*�y1q�Y2�r�U�&b?#6KCz)�.��wf����ͣ�à��M�z��\�@@��ƣ�S��*��|^x��[6�8V�q�"� kA<����u�6ƞY��C���h|���+q\�P"��/����ٞ������*Ӻ�9��eM!4��� ��=9E03 ��#_/7��z�Nx�iB㻌�}H_�8��<��X8�>Q|�7c~r�|C�)�m�B��4�+�
��s�1晼�U4��'��~��dg q?,�l�;�b�J�ϓ�#l�z�Kk�� *��D4�<R��&�����.��'���6�8�}rg�W�g�W0�l��M:�ށũ5�F����\�LF�R�J�i��b	�%p�lY�en��1�L��e{�Ѣ�S �)냈�z��76�v��nH���z��U��n�R-'��O�NޕV0��o��X����jE�Pd���v��{���V�R �J���)R`��F���ze�T���dUǑ�P�>[��iBl�91xC�F�7���j�!-���3���e{q� �׹�#x&�r1��R�g��3�Q_�{����P���:I�3p=�0�Φ$r:m��Ƭm�t�"�`Y�.����)��G��D7��#�U���� <	��6N����RjUu��fRFZh^��v^�i�M�͎n.��~��n<�jٕ�6��@�@N�CC3��m�_=�iKQ����36�Nʞ��~e[��H��-)b�9� @}H&%��PLj����#�p23C4uPWZ�����s9� ���nWc�uD�A��8Xj�lC���=%�2-�;	�"��)�F��Y����:��5���[mq��.��)Qst���FC����͞�yc�ڐݕ�)m(���;k�Zب5n{����7�"�̈J����bU���
l�(���L��$�iW=�fM��+'��6�8(�
��D΋B��g:�ή�j���R�� ��#�%�k%F"�L����� 5��GN��@���2�3��v�o�3i�C��]���n��ھjh�L�ҨA�Z�X��|u����QR�l��b�����A��|���5�{�;�D��}��Z�=�f/���t3�y���޺�2a��0,��99;�W�`��+��^3������=^ڭlu�S��fs��$MGK�P��a �j�%���t����ln܉d���F��ŝ����\.��q�ā��.ɻ�ZZ�F���.�J�j���}ix!6V6�a��`�;D��%�
��$s1��m�~�<Ҹ�j�^��;/oW��q��7/*�)ȉ����O����'�u����L�#���t�6���ƫ�g� ,��P�1��0�+���JĆc$�����pMIK�ǆ���C9%���<Y3��[ŘLK��Iq``0�S��g_�J��F5���/�܀δ�>�Ȍ�~�۽����Ԁ�n��h��;��<VD#BVܰJ��K/�:���������X��@���S�!��.��e�
�'Q�$�h�n
b��8�fǶ���ηZs"���t��t++�o٠��-`,�pKpD�BD/ކ/�/&n����!�x��g�ՙ��<�p�g897o�f,����52v�C�2c_}?H�7r��H��@��\g������k�������؀�K�g�` �|;�~t�2���F��?x0��t�|�����1)�O�������1ࢲal:6ӌ�<EY٩5kC1� N���%'i���P-+��������Vd	�(����p���؟J������
 H۫I	��]�������	�ѵ�Ḑ.(��_5�������̽�7��"�n;��&�ݸ�|��c�1�٥,wj�<�esw�ӝ<�K����I�aD��|I�^���2�İ�k��7����$��)4v?e����>yc8�MD�S�6Y+�h�='�@���#V�I����b����qh2�{Y�c�'���(
3Ć�B���'��+�D��g�f�GP�1�#�6�X�{�@3�F�ݚ�5����wK�&pJ��n�Q/��� P�z3^aQ�:�+U.��h��#:�,K�Z
����8�/@��S�>˼��Л�Ú\��V��d�^Q�/�xޙ��D��޾bv��s���V���"hþ��[3!о;B�q����Dg"�k�¿��8��Fy�C��Lzaf�NU�lsJ
�3�*�n)6�HxP�4 ]����B�ጞ�A��ke��@���a邟�æ��E/�d��v�U�4�d���V 0����o���E÷n�T��������.I�z"��\a�H���)�֠�v�*e.(1[����	}�ټ����u-�>(�B_���.����/&oMH����
,#�4`�aU�Ptwu^v���[�m�

ҿ�͈�7���@i��o|7Ї��_uS
��x}�gi����]�����Nc����|<�?���!J�BEY�m��*13�՛@�zVm!1Q�xd���_ZG�)m��2 x�KC�\r����s+h�F w��X���n�3�s�2F��(���;� ����/3�
�Hf)�	�J�]%/n�� q��T`������-�1�4��f��!Fk�$O˭f�lxuZ� �7��>�δ�<�B��t8Zf)y��'EW%?k��,��H��_��3��/H����\_���d�Mt;%�7�|�k���� �����`m켱�hA�κڴ�b�{�:���S{���Y�	M ��Nw�q'-՗�����^�d�3gǮ*0�Q�!����U�y��/TzM�R�Ȣ���N�}x��+��K�N<�1g1�lQ՜"F�j���a���?��t�2���5��X/�@D�If�`�\*�X��`��r��Lp�	�^Ñ}V������PO�=ۚ�,�`i��,�����K9�l&{�v�4_����?�xRX��ح*���H^:���(DJgN�磼�Ӯ��29}�vXE����"�҉����!���3/G2:� �O��i��_9��q	���EJ��#��p���N�^��O�"Aay���N�ե�cSE���Q���4C�M��.���x医�]�d�P5n�xʎ�s�,�S|x���/�g�T2�Ѕ��!:-n`�2����U
@�y/�ef�}����F(r�_D�E�+�5߽\F��j�k3�m������&�����@�|8���E̓1�Ƣ���s��G[.��ِ��3@�/bWA�}��B��Ԍ��pY�*k��O��e���̗���[�+.>I!�T�Sl#�ˏғ�G��H�n�b�^;�<L'Qra<��w�Y�M��S_?��)��R��~�.6)�& ����l�di�ј�w��� dBh��������2�98��eŲ��}�5gA����W��kI4|�a�N��k��=�ߌ�7�9`��,��a�ڲ��A��݂q�`f�K��?�A���A�-�5�.D}dZ|jQ������	R[���X,ΦW�BTT"D�}�|����9jso�)�ls�	^<�h��4��4��-i��jS��Q$`��Zeg���$̴m�R�A�@a����
�֋8j��u`g5d,D����O�@�ЯHk����4��""�����_2��v�d�]lu��i�5��� �P~�
:D45��a��+�%���΁�i���^*�������o�c��/Z�%'��*a �ddsN��Y>���)#|X����2��Sw֓~�c,E�^����f�j�FR�=/z�>��O�k �f��bړ8�9�쁎	Ҝ��u�P"�������b�Vpo$h������ �;%?���K�ak��o� Wo$�䂰p��-��=�g7��j��n�Q[&sTXx����[q���9)����IJ�V9���TL�3����:^��������a���q���²R��{�:��5,#�?��g��j�+���HO��E'�ݸ��`�o��md2���Q"�cvU}���+J���� �pҗ�{po_�[�2��iF������c�'ݵ#վ�:�.DH ��a���[�7��rO~oл=D9����FQ_7��L7	�G:�@�Ⱥnp�&�s�@���V����dr0Yߘ�M�RëV�0'{n��+�6�^&Wf�)�dk�$,�ӿ#���q��K�g( Y��R@r��+Y�N1/ )v��8��r�����m���2��o�:����
 |5@���5/l�W<��Ч5�A�i����&�ك��?�(����*�h�o��&��}^�9���,�$�[�G�L�(+�[����*k�,����P?ke'#NmV~�#jF�~!õ��A�����ti�����
���)��d���A��O#7j.g�0�������w����L�$�O����ږ���פ�E�UZ�	�_��oB��b t�ZVS�7�Kh����[�7;����ӭ�W[X��d�s��>oG�M몰zr�x�&�����ZÉj��K鿟b�HI���;�9��Ց��G��Ph��4H�J���]M�E��ǟ�mع�ۺ�¯L��JX�������`��z��{�^��s�Ȧ�sF(���Ă�3�����'9�r��)�|���L�>7���;�G�ͽ�o��И�C�!NB��Uh��`�/�X�%l���y����B�Y@;����!�����3���. (w�L���x󋰼k><<��,� �Kb��/JWU��Pjag��d.6� �z+�/yX�o�өXK:d��,�!�݅�z��m9�%�`0)�K��_c֚.fd��
����eL I�h<� :�X��D�{�N2��fl���LC���L��ī���<!��+����9>~z�0�?}b[���[���np�'Q�u ��L�[5�F�Y*������P'�|���W"�̜��B_����E:���!p&�!�B��ny��Cg�p��mW�*�X8�@�n]���p��#M_��m����3Sxt˾j#�E�k#Ȍ13�ˇ'>���Δ��7�]���1)