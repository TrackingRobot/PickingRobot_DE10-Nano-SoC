��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�������+�%ix��;��-���y��6XM�F���
]8.�"y5��[S��I~o03�v�4�W�����x���W��>!�3�i�/�T���Q\�^u���?��bU�I0�k�Y��"	���Y���n�I{�N�Y�rYntf^t�^=���t�{[�l<hX?ۯ��R�!A�cvE4�A��|��ی���1��V�_V�k�Qh����==%�BncC5-}I�J�^�t)H�/����
�����J����}ȍ�N�c�#H�6?�7���2b�����Y"D���B�W�V����.jq������j$]U��b�}w�FG�9 cR=��"sOqWW��ZV��1���9M�QR,�#h�e#ʱ���]#h���Yx|�{/n�M����.�+���c�%����4[o
��׍�A���mW�8g8�F��R�-3T�����)AQV�)T�4�������L��Al���U`o�X�xԵם/r;�9|xv�u��G �����#��;��݃�j�ا;�JH5cy9_�����*94�����ɡ��7�*���x0]E541���}�;L{x�a������e��|���E_:dK7㽨Ѹ2�͉���&����+���j�����HY��NQ3��g��C�b.�Cَ��y{�)���������?_��g��B���S�+�!���ᚥR��%��*��θ�� !�bۇ�����!U
�R���>)ʩ�7���.o[?���\&-�;���F"iz^���4҃�&م�c+�S��"����q��p2�lN���m�j�*�2mn��M��z���u�6�I+�c�%�jf⧦¢��W��WYȟAٌ+E���r\@�+A�>�<;��=G���mM�QȚ�/�1��#����K�����S��/ɵc���x��wo���'i	B�$��S�\-�ހ�Ď&
�N�R��`L0`�E-�x*ð���o,
�DϾ�J9Nb�^�I�)&"�;q���&L� ���R~o�V~<2�,�H�̑^7p����~�L�BTw��	�=n��dS�Ȭ<S]����Ww	�β���]���X��Q=z���S�(I�M9���i���n�����!v�W?q�[�T2�9�
�4�n���sLVǅ��a���Z�w���\Z�F�,(T��k��`��T����� �eJ�9�$���2�ӗ)6��`�D/��Ʋ�N���޷��t��0�(�+fE�MR�ɴđI���]K�a�jF�Ԅ�۸/�>%�8?p�\Vz�e�������#��\�M��Cz�,>��o���[���̰��q&Q	�Hx��T"}�|�ǲ!��4[�� �?�|ѭU��xO9��w���3����:���S�����!��j�g��w���9@�o���q�ꎼp�`'�&��N��/q�K��q��3�7�g87`�f=�J�b,B���w�kghï�$�OL���s�ا4?@:A���60�w���9�H~��;�]�I�ֳ�q�S�OJp��U������;�>�����'�@�"��'���1k��;������±9cV��g.Ʊ�?" �eӲ�<�=�jK0����&:z�[���,�@�� Iߟ��"���R��2,��-<$����o���iY�F5�%�&�Z���o$ѹN�(pBE �?z2J���%�b�cpGn�rF����ӿ���Ρ8wC�����)k/�����6���J/[�}g��q@���M'����p����8����\ ��p�ZM�g�H�������U?Y�h�C��{D���@]��_, ��zB���i_��chE�y�kMه �;*��QF�����@~ej�=�����C��C�ڰ`C0LH�\8)�������c�(��d��QԴ<�t�(���`���NOsڊ���8
m^q_iJ\�Dȳj�bJީ4�ZԮ M>���{�����|VXӊ0;�Ea�< �+h�Y�v��HӋ=E�t�ڽ+��~@�Yگ��c���%�a�38&5���]���ܔ;"��3��@��Q;�Ӳ�����_)hʥҝ�9=�N��S��9ǽ��_5��q#�C�?��)�a=Pn{0/��Y�n��'�S̗�v�Y�r����l�>W-b��*b��l���֨}!��z7!m�+�v��3\��.
���Y��.�φ5|�G?�3�{���/�e��Q�d��y��zN��L���UB�1�D7�fJ]�Z�[w`v�*w��#�i3U�pM�>K��W���1���i�Ȫ��2c�c�g��[,���K�.l��4eQ_��>PZ�B[���rQ�ia���c�O���3P
¦>>
4M��84���(�x�;��]> ���~'&�2�^�
���CB���`F�МU�WRBq?: �v��F|αŁ�v�䚻)hO���"¨#V�Y	2r�:���j္Y�����9B�jS�Ԁm�=U�B�O�K�=��+	A%�t)|��~Mr�����7T|�Zn]ƃJ�
�f��I��<�⪸���㞧E��/��x���.�%g"^}�u�
�cbDJ2�f��T��{��:b�
+�L�g�i�N�fB,�C($��J]�i\�s����.��.0�c�b�=�I�>
�����'�� mv��GԘ��υ�CR�r��P�t��������p_����o��8I�rq�k+=W�"`�+�2KK<gۏ���.��G\XP䂥峫�)�Fa�K}����fd�w����a,8��e}��<�>�qp�Y
���݄�C�Q!S��K8��Z�3�~�g��� v�(�(��<� �c1�Y��u��
�k*' ������%&�رz�ex��╩�[͇qK7Ԛc̣��@�72�v���!��k�����m.��G�:��F�u������'�]���oE�m��c�^Ḳ�7����|�}I�6�
�VV/� ~X����_�X���٦�A�u&�8��6�ϯ��>����@IR��;��҅��3����F*�%���Ɲ�g���vx�o	pC����;�0F(�U?5���GpD[����P=��+Z�����$T�b���^����Ѹx# �b��<;}�=U~�X8�e�J�oJ�Z�z�Ä��t6���D)<7�$���vt�ᒂ���U�������]/�N8��*{�X���s\7.��]<����ۮIPu�l��q�,�9S�*�W|Ny��4��݁���x�xV�c�|�"0����Դ�q&�,�a���>���}�ɲ}�����0�)�s� ��N6Dx��wЍ1���B��o�tMS��N{��E2ܗ��y�1M}�T�5���PU[o�4����>���|��݉π���f%��C��0������Q��!(c��N�S�Pܒ��:��E���MF1�A �i4������������_=tWC����5�k��QYa���?N�♒&@r/zWQ.�@p�:��x9}I�� ���T�@��8��A?:�o𴄮O �˛��C����Yx�Rg}	�@O�;�q��kk�Y����(i@׭A�a��qpg�MafU�T.gy/^`�q��S?�	�q�u����Ė
5+�g�@ph��
z��m6�B���*���Wx3�ۥ�QE�*z(F#߼�Ƶ8���Q�Ae4�.�? @T\XN#�XM�#�SǂI-b���Wo"��U���XO�~�tC%�AE��t)��%W̲�0�z�S�[xG��3\j󺨄ڴ�QF��m���\L�'e��~m��0w���q��/�0P��Q��Ͳs�@�?�:i��0yY��}��*ƻ��R
���B�0�F>%{M-�1��od4b�MH�9_�7\~�thie���A�PF@�i�l��T�Ľ�s9��V/(��jP@��_�6�]C�M����`�\!d�������$��SZu�"1��hr^Yr1[���)�!��;�UU2=6Ea���E��o��]�!�Z�X�{wP�q�ԏ��q�|�כ߬n�T�˨���)q��$�NȞN5Re�3��>�?K8��:!������:-/y�8"I��qr�
X������B��ca�s|�M�����Ýw��h;ˇ/�4��ì����:֍��,�ٟ+:����Pt[`�5	�f�-"�_�l����>��ͼ_0�axw���f}��>���5}�W``��fkh��If�˄3@��U�g*�]�0Ab+LFP�H[���b����K۵��W��P�w
�*��s��ѳ����=j�ΈDuXZ�\���'��T������'��x:�BӲpV��{�,�r�=�r�����U�7�)m4M�G�=�)��LQG���Ĝg�Όh)7�������P��Q��+9����PO�/�e���.�e+����}���}�ӽY�T��M ��R(�+���MB��`d@�{?L���;�	�"�c-�I?�>�J��@��Z�V��;�QO�t��Ӕ�z�?.�]���\��y&�1mG�2�W�,f`�����~��A( `�*ȶB��|�w䘙����d���;ʪ�g'���n=V)Yp�Q�^xa|s�]b�1p���ޤh�.��KZ�����«���A6%��m%��e�]C뵯���Y������Wl��|�`1"��+�/<Gd��oM�0G�+φ�@���{'��tRW;��%�k�=ѝ��R��/\^� _c�葮�����C8a�g�6��Nl�֪dfۂN��d��iZa��r���&rS�Oo�9z�X0<Z����x��������2X�FΆXf����&k�F�͎���Ԕ$G�9�����cm���Ƕ���7�������P���H�?�����^:�i(]���O�]��ea���>谓2��nN֥�w�����ԕ:r�K��V�u�Qlq��0Ţ��WL���̓��J7w���=%��0��'� t�+9n�P�ث��%@�cR����Z�[;eL�a��Xo6\��&$G��q�܋.W���s����|�t���kŲ�So]���9����	��=����
���^����6)���m��t�\�QHD�W]&%�����c®��������F�3�S/��C�8��NJG����Q�����-`M�TX�rg@��̍[aոˉ!l��}!��y���b����M���.�����P	�b8CN]N\ǒ�GL'�/Z�������$���
,.�]�C`w�2iWa�0l����e�X����m�Q���zX=쀿�<���G$\ߏ� k���8<�n<f8+�;$��p�->���Yy�
����}@���k+���&~�7T���q?�Qg!�m�O�j��P�}���vL�iQ80�q�����ڡqQ�h���L���A5ƭHu�r��q�	����i?T+����v��ձ��d�H �#u��ڏX��p��e��s�^�90 �&�;ܝB�R��Ӫ�j.�Ԏb��F{kI���A�+!h�.Ï�۵�2�-�Db�d��Z�=�"<·S���U�b+���h�2I��a@f�g��)�S�=\F�h5�����[�\9�y0N��!�;�}
y�`]
yS	gG
}����;�i���۪g���T����t�3R9ç�E�,�OF@;����CRs��%��M.nM�d�R�q���q��}s�u�R5>����ڲ`����b�W�����BS:Гg@[>����lw�����!{�E_dH�~oMS�KH��"���b����|tNAGО-z~�j�`��&�X��S�|��Έ?�@���Dm~`��$���i���w��⎑�d�=~�jr".`�j�޸�������0����=RR��N�%x���h~����2�5�s�cC��c�S�
{�؎�27V�lL��~�Ԫ�����jY<�fD��2*1��C��SY�p�K��F�� 3޹�7��.��G��M�N�v�6���*��g>��,ԭ�>�5�QP�7_��.��&z��L�(�A�Y����%�(��} Op�� DF[��WN�MU��8rs��ʬM�?;K�:jb�orc�~G��Ү�}�����٬/�㳺����]` 	�+ؖ~_�<�П a���AV|�
-���q�;-�TR6/za�+�U�]�g��D2����c.<wjBϞ^ܪP�ߚ#r;�YW�E�3Y�Y�.�����t
�����d@�ůt%������8/7j�%�&��R{�qU�@}ь��6<�7Y����ǡ�Q��� ��S&�&����_A]:����pl��!������h��h|ijǗ)�.b�3X��E��0z�'�E�p�=7d���	�.<L���v����cTg�yl�(Ӫ�y�j_�&H��Gg��@/��m�>ݒ�l��V���P�K}k�0�{�@y�d�\�^gk�8C�|�~�2�k|u���E��J��EA�n�rT��˅ڱ��^ֵ��u2�/Q�ՒTv�N��3aF�ہ�]J�٦�!����]ar�N����?��'�:���!n�aN��ꂞ��Q�*,3,���*g6�g�ʌ�9�뽱�TJ����<�i(�-���Ն�c��O�%g�q&�T|��0���o���Nv��2d�a��{���1/n1�_b����_�`�:��7ş��˿m���.܏���w�c���H7��_�ɮ{Z|H)�Q��(,G1t	��4��K8[���O<dl\R>����h]�hF����v��׍�A��Ĝ`��v�bl�6��;�����_V�j��5�W>F�2O@���y�����b���	po�;�����TE�J�H%�XJ��U���nN���e� ����5���+�f�歬���5��3��]��]e�o�O���L�Z�lM�25�B[yi���iJO=sɄ��`�n��~i��
�T+)nYpg3F���k�v�J̿N�\��0A��$�����d*3�%ێ>�o����,Z'��N��B��1��f�r8ڤ��q�{+	���s ��r� a8�aE'̿!�j3�Q[l��Vy,�wX��M�_u|�&��ͪIjq2v���Oi�	*oh.}�o�5�d�2&�`�(ǔ�*�U���r�7ĸN�<!�+_�V�����>���]��=�{_�����L�9�A�G����뛙���',���>��P�����'��C??U�����K�:g�$�8+7$d����;+���������N�5�2p��� &� 1ND���d��w�s���v�|P��خ���c�����J��%0�y[�n�-�^)�j�D��,�@�o�@�;�[�v�{���j'F�[�l���b�H^���R}µ�c������"�ٷ�LV����O]�$P�MZ�k�,�H��� �O t98?�b����u|�� X]H��Ƞ��ވm��C�4��(x����0y�	�����c> ��{�wm��j����ECa�?�x�aB�.Vr�y�B��u���(����sɊ^F�����N�1�m��5�2(9�Eһ�դ >n���2��<�cH��9��J;��C!1��Yѥ����)�q�-�<JՏ�a�
?�2ڕ�j���:#�������&���Jg�u����x}�h�#�dW'M�L,�{����j$�_C)�8���+$���\A9�t�l����c�� �2�j�	r�۫ BFʺ�K�6
�x�I��[�(`�R.�{�������h�_�nP����c�Q�>*�N���WӷC�_j����!�t$e��{Z��\V�ۼ ޚ;�/�1"?���ʝ<w�ʫ�ǹ��T)�EP�v�0�~�+�u�`���;��&5a��x��=����X��M�6ջ]3\0)+�\��>����pRbܴ��v����|�W��k�E`�6~�3�B��1L��Y):��tnm)�0��A���W���1�(�8�9�G�ͫ����Ö` m��&�"���p�K�/�n��#{����#�~�Gg"]Jܣ�	�ʵ�������5$P�(U�,���u"���9�X[�F}Fy�/s+yN*�S5�̭OaY����fi����	B�ik�Y�j���YsE7�;�д������R>��!UP��G�ܓ�����o}���$�
N�3�U�������2�*�J$��5�s]�Ty�0(�q�,D��Ţ�0WdB���@�#��^A��p�}�}��,�҅Y�s~�Dqx�<���O�c�><��)�җ.d����|٧�:��B�����슘+Q�6�9��/�8WL���Îx����~ٚq�c�����d�ẹ3R���#o������Z�U��h2��HA�̗�9�`���U����#{!e࿃NPx�*'��[P*�H�z�2B�Hl����w�+��.�Ȋ�#���锂/L���:Af�uY$� �>�ycѨw�,�̻�-�a���<� �h1���.&8,V�|��{�M�����M���捞�;J�0���c9�Y����S���M]GW���j�_-ҁ2�V7���!��R���z`U����\U~{�9����y��(���?��M���P��#��� SR�-�4s�q�p�q�Ǡ�On�a2"߯b$!���:�(��l����|�b��Z&	
-�r��Q��~�J�h ��F���εZ0�Ux�3��"|l^I+�S{!v�
�搊�G�R�~�%�7s{v�m��U�=��d7C���S�V�<��ɀ���X�xF�B�1�E��]w0�&�U͂���*�����I3~	��֕rP�]ӝtH�AT�)�Kj*�'~��U/��ݯ���� �Р�3��(U~��tǦv�%g�ܕ��I���]e����4�)�$K�C�����b����>�@���B��jS����i���t)*k+�i��C���Ϝ/z/EG��۳q��?���ny�=�M�k���w�zm^�Zv���[�LY��	�L�ᓵ����+l�5��~ A@���a7Y��dl��q��[o�乜���:B���p�����ʠ4s�o�]3f���0��1��\
EC�l��v�$��L/�p�R0�'����(�F��-6�V9��"2��[!��g�&p�}$�*K��aӥ�CD]qq��gr��?��S�X[��=!��NJ=�L6�5�,=��{����
�fml�n�fZF('��|��8�uђX���ȩ�
��Fn����Of�uGy��v�rc8%:��QzsF��65Z�6W@vm-�乥�^p�c�j3��@�E)�ToF:Kn����/tһ�"SmQ4��0�2�q��Q���;��%i?H��m� ٻ�(��2�����>�&2D�����(*�XX��6�.6k�2��m������sr%,�V�(r8`�L8��L��b�"��<�]�%.GbJ��t��?כ)A[�p�g�<*�k^���.����<���@Z�-+?re�%�zyV�/Z:[;�M��.C� ����ۂgc�%��Xw�#|�����֤M���k���Einߣ����P��OKҹ0쨾��� ���#3�Y�Mm���?0��vRχ�Rb �����Ź:\�g4?�&B`��M�b�WɌ��"]��%��*�1����\5�iv�f�TmJ�����oTZ��.c�i@`&[TT���̗a��mA����NƤq)�D�Dq,�oh>%U��]'�'��)P2���J<a�^@�zX<s����Fx��%k_��@F�a˹c�j+_C��O���3�V}����J��=���*_�P��"x�#����b���9{
ڪw`�wp�^/=g�H�o��C
q+3t�̓��_~��b~�vH��oMb�����N��0���R���QR���[U�3��_��`^��G��"�YE��&@/$M�;���x��e��<���!5d�W�\!}�{���{��̎g Tcu���dD}}���#F�N�Y�j�ެa��:�����h�̮E{�`�ޮ�X-�'�dQ��l���O"��oR6�q�y����m�Ǩ��~P����ֽ{�����Xt�ߌ���\�ac��.�ur�<γ7�)�H���Ӑ-'x���	��7s(��~��sd������g�/j�w��$j'��EnT�����#�!�}���R�@BŖ[qs���v���8���c��n� ^6���!b�ڍ#,mٽޛ�:�b$8O~�r�?��8RAw����8�\�g�A�ݚ
�qX�~`��Y�YT�!`7_���M8W���� �3��H�;g���4���I�V����އ[���)�^��;^��g��f�J� �v�Jc���� �]$ڴ�.���XX��u��o�f"O�C/��i�5�kK[D��8ī�"iP�f�?�H���MV0�A��rT� 	m.��w��P��~w�@�t���\���X��g�02St���G��9B��K΋�ז*�~<�b��o��@�Y�/`��F�1km�9��q���0ׁ���ߵ�(��W b#+�\Xb�>.��٥'��V���Y�I����[I&QRA�����Ԛ��� � �5$1�ɃF���`���L�($����Q�j���5�Ar�ѵ��1GH���0�G0����:Ȓ�s�;T��Ԇ!'T���[�o�g�(�{L9��[�-��Qfp�d�p7ӌ�D�O_����u
=��D�˾"�y�
�x�ӓN¨���QH�V
�aV�Bv-br�� ۫���$�xF�u�o����Jm�n&f]L:���uG�=@�x^��?#�b=����+g�0m(�;�)�;���/��c��k�s�~�V�S��}�%��1�X�L)�q� ��;Dt��R��S�w'L]	�`Ҥ��1Vk�)�b�L�pȈ��2p�_s�Z�KVG�lP�: ��	�Ŗ�Ѐx=�_�ӹ�(7�ڍd�ٿ�����N�aC`��Ϝ��3��ŻI���	�����#w�O��V��y��>�	�>���͎N?
+�ŀWb�c��Àh���q�y�b� �N��(���.�?�g��7���4� ��q�Ϡ˩��ܥ������&2 ��ju3�1��d}���o7,�C����ξ��xX��u����h����A)��=����fMs+a���ByvM�ON:*Up��rY�����'��0��J�*/�x��zd��X|^�p����t��r�t�R����C�S��I��G�9L�pLF�G�-���)�ۢT6G�'H��&�g
Q�!}ܪ�x����WlB��+���$�x2��s���~�fo9�r��ԭ^%1=xc\�ӵ<,'��]��{jĩM=Y����P��V��E�u�C�_F4[�,V���n�vv�5��1�+�՜ʛ�:�����"���q<��˹�B~xJ]Ω��+d�/�٪Q_@b�FM���\R�} �(!��D���5��v돫��A%�ߜ��u�I�-�A1]p�%���!���>�_/�S�L�>5qj� �|inE�g+5�uV����Pʉs0(��?!Q8�H�_��/��&�׵t T/"�-e�Y���WL��ո�m�G�7�"��{1��4�.�==��,�]�U�L0���#)�v-O_s#u��1�X�D5�_�PkF��9�'���U��'��E�h����"�׸�ä[73*&Z�:�3U���ҩ��7iZo��*�q��F
Ƙ׆���̤n�<~	.���pAX�A.���	�-�5���z5ZE�bkL
�����Ym��[�N�m�sD�߃��~�@rO�A��^�����m�f�ꁫ��-?���CBaݽ��z�O�-�j�c�EWf�ɏ�V�:x�s�S��	M�x͠]7�r�/���lP鋣Jj��ǿs�-�I"��X���_��?��v�q�ҿ���Sn�dd!����Kܖ#�qH�r�q�d��)�gMh��ݐ��W~�:�pry�$�\¡�X3Tkk�l:������ї|P�k��_�����ʗ��a�5h�MJ�����cj���^��c�9_yW/%ڊ�5��НDK]���2����f���eY�7^k�i�b81{g<���Y�a�g`aO���H��i���FV���q���O�j�x/���;_�9
��G��j��]�đLD��]c���2�F��dU����4��p��B�Z<�6����[ȼ��*Ib%���o�oXף�5�Z82f��.�Mñkߖy��qh�F�ݻ�q��y���*nMi��.�dF���m,�K�D]�&P��
y������B0=E��yeC(��!'���¤�
�+�� w��W�S����sV[��z�1����"�#Gn��>>SH� �Hڗs�� =KՐ��F���������S-'h�m(/𛈱�������+��9x���	�p�06��V�a��}/d眇� ��%�{�}�G[�c���21�w��A��p-+g�Ku��R�`���q���Y� M� ��M�� A�2m�Y;�v%���1
]@x�
�P{�� B%�̃�,H����~x����;���x)����6� �nJ�-���@$԰���x^�\�|}��J&�F](A?|J��
�������� ��>��?e�\my�"��I�ϟ^�Zu��4F��Z��#ēM����I$�������I:*C_Uz5�T�y��s�+�������������2�R�ރFb��_�2����?��qX���/�y�� n���wq�M�_����B���Ց'nl�K���(����$��_i�,� �!�<5ݺz���-X��FL	,s5�5DLi��I�Ϸ��D�0,OW zW��#� ��dLUE_ �z�a����� ��v��	� �m������a�OE\Ӕ238��W)�9.����q@��V9n��#��4]d��ӇJ+Ԝ���O\Oqqn1��cq�=g�/�S��i�o�Z8~c�����Ȁɹ0�Б�a7�,n��&\P��$��/d9O�$�S]� x���\��$��w�h�)�oaW�3�v��!b�I7�#)	<������\]?	�P+���I���a���XdA����"'��Y3�I��X�x�$��5��T5��!�-� ��g��H�G'�6��f�̏�Fۛ����'8�����Mc�sb�JY�o�:�ڞ��D�&��>�:h}�ሿx�����}����/��E�C�@sx34ZԀZ@q;}m�y|��#)`$�i7e�����6u0����c�ke�kJ>l~%��V�$��s��ɠ�l�iw�VCQ����1�@�*b��1��*�Q�`[��=�`|	�f[�>��wZ��	L͈ γ0�9z�[`�X
bƗ�e�R0䘆d+��2).6R��Ag1����y��y#0���pJL:�A�;	��1�m��1�}u�=����v�Q`o*�r�p��!�{��Wr�f���S9�(�TI;�����WI���z�9~wɃ-`\)�2��6"@�=w�))j��r=LO�(�>��-�h!A�m�o�"�̈�bY����s�B�V�	JC
���6���-���2�h+��pi7�&K�,��}�b��1K7T\��79,�L}S���J#�B[����Å&_��{�9m��@�,����&[-K7Ɯv�<�����X��i�a�χ�Q��+I0870�<o����ַu�}�A|?�($�5s�J�Ͳnע�+�hpW��D�ef1��m�u�0L�%��E7��DI���!8���,V����n�T�]é��ւ@�w��N h�#*�JIԞ|\���(�G��
W�AfrላѼi[�0����/��:�?ۖ��c������
��>�?�Ng��2����]Q���+P�2>�$�B���Kz$1���2/A����L>R8��K�#4P8Ge{. ��fI�YJ1 �5�_�:6a���"�(3��f����K+;b)�Q��(�X�D#4�θݒ��y����Ke�G(zCZV�8�+��5&��Sj�Q5�@t�%�B,�ч���1;���H�.Cu��ak�EU��йr~q��sL�N��Кmozf��N��n�5gz�B�8��{+h��)N�����#=t�.%K�9����Ň�bFޛ�.W�V�$��Z�!t���/�y�N��?�\�4�CȪ1:d�:ߐ�o�4Jk	>4c�A�N�F�%�kGr��l��Y�����G}��޴0s���4�-d�-����5�c�:����<�P��:/��nPL���4�O,��!~��l����B3>^��.eĻ��زp��������Ed���xx�K�Ug����������zOXB0B|�Sw6��B�bT�!���\xf��^�1�B\ہ�����Ow��v�B�uFP�����#V㺑�Q3��}+ُ`�
���i�tvWVU�f>?y;�.��g~G��qG@�'$����W�"��KK�?~�45�D�����O�Uv�)O�ī0�k�Y�����ף��~�g�G����bI��Z.��Y_����3J��=�%:�����ŏ+�hx3��>�4���i�~\���G��������l�Ŭ��r),$}6h۬Dt6��S�Wʕd�;�ͽ/��J3�!ej�a��[����"�x��ْI��L��9�o�q������r�b�]Y��^�g�H�L�'hĈ�Zf�i�|���r.���].%@���Hz)�7�%�6-�4�6�<�-�Y�EՇS�|��Lm8��J��ko��g`*SC�VՄ6"��� ��u@?��ic�DN�����o���v�,T۳����2S*���s���	a�9�+����������Hk�y� K{j����
u�*d�6�zb�n���
:#a���F���[9|�>��;`敋��pom�e�x_�GT%�ӫ�s�w���釹�T��Ƥ	�)�k�/���e� w��8��,i�8|D �D�6]��%M>���	��I^�]I62�Ą��>���2 ��;b
,3�8H��i߂v/�ѱL�G'��\Apv���K����ek]��}*��X��x����άS�&]�7�i���=�_�s��L=J��l=�<W-�#\z����}� t'�$�A2��f��Q�d�#�8�ɚ[�U��Γ�Z��o�|B�"ܐ�%^�����ƻć�뤁^�5%��B�i�������#Um�hfEW�!��t�Z�����o������̨ҥ��|�^���n�^e���ZmS���8����iO{�L�}W��[�>%��\Zʁ���'����: Վ?a���	�ܾiH��"���P�E�?�����J�keW�����~�����s�Qkw�x(�~@� �s����6�~̰�U�{�gc�x$�g�	 XSU�$&�i��ӳ �u��_��N|<�ه���t�&v������!
7�8�8>hY�e���-���<v"��=�����a�֐jq,L'V�5����ћ�����R�[P���N�:�CK<���������R�����K��ȕh� '��~!kn��V+Y�Y`��7��������^3����3�ćBw2+.��M��6��m�j	$�^��o��G���ig��b�J��̈́�_v�W�_������-]=#M|�v:90K�ƚ����'ع/���J�=dKшx��葰�M�i誩�J������j��o�؟� ���3�L+�]T[��j���;�h��u8��uS`ٲ'٘�X���']'�هD�Jf��;NO+-;�n������`�`Ц	}� !F~�"=����jX�_�ݿ��Q��4����"M_ڝ}���Wdg�t�q�Gj�ƙ4��a��u�]���VHq���Փ9T�F��Tjs9�b�őH8&��A��J|�Z�Z]9���c\�b ��v� �Л�$�pl-� A��Ƀtr�X��P�5j�o���3����限��z!}�o�R�9�K}9��*wE���#��V' ��\��K�6����\MكJ�x�iuK��s��+��{r3|v������:ŢC�O�����\���ɫ��������U�>
Dx��_;��%���{^�\n�e]��ׅ��;�i#���#D��C�*�8��`%���p���Zz�V-|@�+K����e���Ǽ|EK�b��B�[7#8G�)ݧ�+���A��O�~�9���)#���*F(6�.K=�6ʢ��/\h��:�����C�e�xI�+:�ig����9�0{�EY�\/��q��cn�?&���[AC�-ט���Ia���T'Jٲ�1ߟKa)b8ȬU�.M�ԷZ��sg]����#<?��'=2rT<!L*����F���N�x^!��-��	�_ *Ń��^��L�.�'���d�c���iw��'�Ƭ���� ��PT��-L\�E�����l��R�Cy���!����������M(��Q���W���D��������_'9b�V\� ��g�}S�#U-����k�DN��i�|ī��#``�S� �Ż�F%m

im�q�joP�[��O���Ya}���ڼ�U"b�t�Cй�jd����X�{O鶺�������<��_a`,ӭ%٭�	y���k,�%Ĳ��)�o�b ��(gqi�w׏��p���X�*r�5s�i��.�߇��x�3�j��u�M�`�k2��nն��w����L���*����9y�&���I�l�E�rf��?SZ@X��#`�'E���)&�*1�I��`}k5��t���3��,�4H�M���s�ʙ���$9��$�~[��%Pͽ���Tw~,�U�L���'�l�z�w\G�S�(rkn$B~NF�o��������93�����>k�9�y�[��:P��g�$��u��¬5f4�,�8��{�K[��t%0��bV�a�����I����F�Y^D�LT�4����aM3�R9d|OJ~	9���#ɪɠ�i�ߔ�Q�V�7��ߐ�3%M��w)$h�)�N��N_a�9d�\. �J�ms2�o�/0��H�����+Q�Ο}�.�Z-Dƒ}�v��E�6<Q�\q3�t���E�	��i]xL)t P�s���vz}k��E�oyb��}�	��9j3���3]��Z�����vy˃b��n2$'^-���9Z�q�Y�����)��+�B��>��[;��R���T<Xn\�Rڔ0Z!)�!5��`�H���"�a;By��p��S��f���G�&�`������/-Bf��?�y�=5���y��*���]��R݅���&��T���� � U���Â:�@-Re*�0�3rkc��Y|=��N;pIRop9ݬW�PW*t����v�t�]��Q#D��WP��$Xπ�.3�������BU,h-"���N�.^�V�b*�'�
�2����2���$#i�9}`������,j(m��<��仆�5��'fd�!C>d��F���v��ᓟ\*V,ļ��rF�n��n���1�kh�?���G��Iv<a ��[��Ӿ����0O����v�IF��aR��G�$"�S��OV�̓�-[uf��%++�J�G��v����	�d��9?�2oK��,��v�b�^�u��'����k�^h)��QǠ�	f3n�4�r��/�Y>=����w��ƴ��s�N�Q��,�@���#�����*9�Gz�U7���:��f0�B�nr����	>H+ӉDT��Z&�U�/�8���7>�(��1�������Q]�_�;��M.�s�9�g����9}����9c?յj
2�%z�Vp΍;�����Г(��&X���Rۄ���*���ۡ	�j�J��Oc�e�0H|T�=����+��m��9�/ظ	 p\z�,�]�5��w!p_a���*��}S�(D�¨o#�R9��g%ß�5�H#�u��w���@C�H� ý�-F�D�4�5@c�f�'�p��6�m��������,Ĉl��Q��+�J���vĄiP�b��7��y�"1e�-�V6c؂SD흶�/]�Sٙ�~4hё62��t���:}0~�Q8��.�9��ګy7��E�(�K�%���:h9��7}���_��x%�q��GB<T�ӥ?j�Š.!ni$���x�'ل�o�֥8QmF�:J%Y�f��<�:U"�n'��O���ُG�t7��exe�>.����A��SH��u�ӗ��V�+uio�!a����P��L�^�,]iT�]0Qߝ C�����n��)�d{s���H��$���w�k ��Y~mC�l\9�0�`�t5d\���6ѧ��u��}{�q`f���d7����1	��κҤ�kj JD>�0�){�F�si��5���r�5���������9o&B?���mO��OD��p�v��7�����+Q�.�1�G���U��c�S� 05��0U<��[WC�S����_���e}�#���R�zE���Į�J�I�M���i(B��ք��^�^ϋ6��5��6�ܺŎ���W�d�>
�q�E�4-��M���Vg��\?fʹ1��C@���g�5����V�d_��`�%����/���� +_�Jy��CF]�@�ޟ�&Mӟ8��s�[ok�>`>���{�Q��y�8LpW��XZZޫ;���g�oo���}J��۔#�"ԉ�sn(��V�NS�wc�E�4%�tSB���s9;�t[�k�x�U��zT�~�ci?O�d9O�%f�Aep�В�G�� ���Y��u��X��*јUs��t4�~� ����o���4�2�"3��"P�3���0{�5\=��g��?
��+h��LA�\y\�Xwzf.2�4�_<�/�os�A	�-��G�7�F��8�7B�@��6^l��h�F6��!�)2��K,��ֽD�*m�ޞ�n�� �Ӧ�u���>9�ͺ�n�ș�ݳL��(a�����neNv�[o9p�D�~@\�_g�Ƹ=���P��>�0���H2�w���|X��w�GL{�i�{a?����hg-��#'�P[r��%�b�"U�������c�mI���FC^Lz�A@@wͶ�w%����7�@�]`{>���;�؄~���I$*<���Vͧ7�����at��VC3��]�B� ��<���m[t��|*:�[؂�[��l�^��"�{&v��+/��7�%t�V R�(��cD�G����2r�u:�Z�K�pI�f��N�C��4��T��T���J-s�R������J��1�x��ן�@��(��PA���Y�?*f�k�%8�5�e�酲*������7�>6�k ������c��}U��C�NIG >}���{�v�_��n�%h��GE�������ce$/��K6x��m��<���i	��
F+�4�T���VG��ͻ������R��J�E���8ݻw�a�G$Tb��u��Ec(< ������%��t�e�^&�ơ�en*+$<Kxb*��jf�<>���8US�'�u�ǒNC_�@��L��Bۇ�$��)� k�O�^/����w��,����~��1�T#\.��8��SΞ��7'�L�=���>�?��QKC���+N���8��C��k���U�z��չ�t�_V�ɨ(�@�Y�M}Y��2��1��}Y�_}+��#��+m�pI�Qn�6�m֞����z2q�m;/M3Ruo +~Đ�~Y�EI~ �t�Bv����F2�4���(	&$����}-lVE�o8�<)�ݥ���B�ͨ3�1�w���U���]d ���E|bK��~�'1��Ll�gD<��i��"9��F�mR��41�uWR����k>6O	t���4���A�c�c�S������<��e�����Z֖�DF}MptS�/	�fK��Ůl@�څ^S����RT��B�P"�I�p�Qt��$�Lv��|��7��6A7�����g20K��#ӗ��)m���$�
��� �x�˫)R��]���u��b�9������\��n��륋aM����M��wa_8G�J��	'p�$.�#��:l�eFǦzJ@'�����H��{�}�G�1�"�v>��'�׶i{L]"�bB�����6�	��?/ @	2��ʌfuw�����O @|����%T��M{� �$�Os^��G��0ɮYѝ��*^�Y��M��]t��w^egO;HC�%��6�t�o=�+!�D�[��E*\0�?ѷ����3<
�s���}!+�;�`�ۃ|���5iP�<'ʂ�U��).k�U�0l�6ipуZ�@� �4��e#��I�::\�ӭ l��t�Vu$ֻi�ѷ�0H=ָ�y��I:3��k��ݔ����AjE�%�g}(��1
�cuE�B��j�>�Õ���W6}:}��Kᩭs����>�P�?)9��}���a�%���ⰲc=�B/Wh��0VP�V���yꅫ�y��O����.��#@\�(߃1�����W.@7�MFL�6�.c(�Ve��:�4=���ǌu�s����iQ��ؓ����v)�ଓR+&U��� �nfP�7l�ݍ/g���fC�^^A+�
�F[�*'Wa��i�ë-{>���s�r��;��3M��9��wz
���ZMq�4d���f�J�3�C��f���|#Z`Bn-<�z�)ڏx���z��nZ�8/H� |+�� v���������q
�E*�������>�G~��aq	F�IHly�š����CN`�>�S�N�$��b%����s�MFt7�ڍ̓�aĨ�Z�W��[��ؗQ�9 ?�yY~��qж6�4;��/���(QD@QH>
���/�J.��{Y9�BX]�D,}Ro�C06���o���1ȹ�&a��+cY�{c�K�Ѩ��_�����9������(zm���-�No.�`=[q����e	��u�B޼���ܙ�[#U hr��]*z�H�<;��O��՟�\S������UM��gj����{���[�V�º<7���ˬ�J���ۃ�_wi��Ԓ�"�<�hLeDV@�C��ѳ���%�O��n�N�2���1�g> 8����-�PH�iO��4����~�i/7����a�SEG�	+dE��j��e6�1A�u�$�2�L�o�ϡÝ���W{�Wkh_�����a�&�4�o�,I�_({x�l0 JmH���8j��@;����{Go��/r�ۼ�m�7�T�3ŲZ^���ꩻ�u��� ��ʃn�W���4|��V~�T39��)��C_�]�؉d4�G�&^���-0xEf���F[�ɤ8�Q�1d[ҭ4��c=�3����\�tڷX,��GZNTy�y�|�L1$xj�Iw�>%�7�g�RO�@h1sdӿ�=�ڬO�|����Pa�6Z6��9_h��[�A�GD�S��ĖB
�0��'�qP�ͣ&���O��������X�����h������=H�M:�ֈQ_ӎ)i�JPLdz���+�����%�bBœ-}K}���w���!�-;��}� ��u:?��>\�\
����SR��*����I	��V\��0�7˃J"�HsК���a���O��M���kВ���P�\4����əB�����d�^^;���h�yp�ӳJ]_eu�Ks6M���[��Ո��
I���t�kӳ�$j�yх;ܰ�褔����ϟ*TC�*&�L�D��4��/��pEX�����lu���v�B���5��)�I_�Ӿ ّ��a�Td	b����.>lZe�)	�Nc9w+]):Ma�ԙ\Ls�fMIŞ��=�HѼ���Sb��{�������	�:�	�+�1�B�M���r0����>���&q�W3V�6 �_Ԫy�J9p`���)%���k<�۝%�c���j'6V͛ߣ���Ԟ$uE�u�Y�8��,�a�iyf�
VɉE	�d����@�y��?� ��wɘ�k�=��W�Q���'D"��ܓ��.1���+�$�j�ֈ�<X���a�m0��j��3X8o�$o�㙋v�v$�=A�-�I��y��9,d
�$1�(������}�ё]���sy�(%�8%tW,x��\����8�Wr�8Rȴ��ɾ�pu-m2���B���Ơ���u��V�8�?G��蛠�~�̱�T`�%�e�t�A���;O�!,/4}�]�߅*'uzsg��u���)-�:JكY���」��?���w��6+@�6���0I��|��'�z� &�q�qo`žef�����X��Gvj:NM	�p�I�Lw�u�Υ�9n�?�/0��2�L#�y,�!5��w��|���W�J�ֹ�ƺ�%���Ro� ��|ϸޙ�-�A8�e�
�MR>��M��u��8(5Bq�稚ah����\��.����C��k�;�րGkC1�}?BFh����B4+Pt�m�����M�6��^;�+3�D�^D�6�s�2��E�:qerL�;ˍ&׎gr61�y�Wx./턶���%�d�|m�	qҔt���Kd���:a�u<v��l��IM'D�J�c��NAi��Ӊs+6�~�{����K�b0�w�V'P,9+8�wŖ�-K^`�P �/2�85|.���n��$چ������B��O�d�~�Q��)3�	��N�Sf���W6H���R��^�l�k�M��\�M�GrI�h፷�ic���W�o0��ٙ�_{�;��{��$��j�Zr�Ш1P����)��mX��~������(�)��q�8aA�x��݋ؼ�@z�k���;6``e� �14֮cy Q�'SF��I����q��ň��/��W(�FKtcc?���`�r��]7�,��~��a_��N;w�Y  ���yR���+9
�w�������$�A�LE����	�AYs"��N�WsUUY<����X0C��Ez~� |V:sn���0�9v:��<�c��T�.��dB'	9�X���W�4[+�
�@�%C����l�P��H���.�J1�	-���M������W��ᡨ�ɗ��ب��SZ_s���-K��M��;5	k��!���KӅ�t�5D�3T�R�1���i���%���U+_�r��@��SM�YIy�F4h~ߗ'W-�6�@���o6%�e�}����8É&��C# ��"����)e��b�V$�$�}mCs��Q�����}�<6j�ר�2��b�������@F��B~���^w/"�@@E�����%��?�"rƻ��*nE�z�PmX~Q�����<�TS�K�����݂����ں)�ǔ��w:����t��6%oI��)9��؎iTڐ	����zqLn���w�P<���Oo�s�Ύ	ג��'A�x%Ѱ�ZE9���g0s��nƗ���8>�F[��J���G��kA.��_�r�w�tv�CXD8��x�p����2��
�&m*��� B�P ��p�}�׈*o�V�2v���	��}
��yR�����r���=�ӹKĸ����^�ؐ7����r�}�tu9���ߨ]��f��榮��u�p��]sX?��L����_�	/��d�=�`~�`��nY�E�4���Q����	m�Y�8\�	Ed 2\��Z=]B6�%%�Q;3g#�O��ܳ)�ک �s�o������ᵮ�Pqx�'�l�m	v�C��ְ�Xr��ej���|�V��n ��)�/�Pkl��J���W;�w���J�c1$t͌���3y��Kj��!�׽g�aJ�B��ڰ��:@�U�3�	r�ƻ79)H�H�$��Mh�/y>c5&�C�W�oo�r��C����:�����x�S�B?x*ݰD���吸a�B�5�b;�R�v��!=e�`�rրG��[,��+cs�/�\��z��^�$�e����9��zd��6WfST�aY�'�U�W瓬���us�͢��+�ʏ�-0ЈH��Y��� �y�;�hG��:	;��^�x�ys�L��٪�󈆞�\��P$u�WĖy����N��P�_u�&@�X���KT��Gh��~����T�/�SsP���4l�>}�U3�"-t�ċ!#S$+��]r��$;�q�('���#��l��C7wc���gTx���k�,]��,)m��X"�i5%{��|h���p��C�k��\�<S��'+���߇yK�ک3�UG��?���^�2��GWo��c���@���:}�Y�,;ZJ���ۺ&1ړ��
A�pT5��}�ɫ=?C����y�ټO[�$I݌�g�;�a�H{�*�~A��G`e�>�T��/jc�׶�����:,�o���R�]>&� "�������W}��_&��iQ�I9jNz}��5'-�SJ��TO�a�T����1N�u�
���%E_v����=?6����4�_�v�> �����w�f���\A AY�|���@�ɳ�.�vi�]5�09 A���R�VTc[d���+"y�Hh�?�_�Pݓ���9�{��'����]���(?Η9v�W'~�j�o�/ߡϮ� ���f��go4 �Qe��w4^v�p��rhkN
r�O�^�`��W�� �Lw�BZ�΂��໻���d뮑���*վ�b����r}�퍭�����!w�Nz��pw|��@�Py�8迁j:! -։�]bW�i ��]Ls`�t?F�M��Ή���k5*D�� �Sr�r(��,iX_�O;8����Ks��=tx&����7�7.�øWCa���2�_ro�O��T�&{Ih0B�M�#�A'��h�"'�;�p�3�8� ��`�I���f�q}��ۄ���L�u�FH������5��v�O� HD�g���[�)w�tX=��΄����?\Ҫ����@�d������1�W����#�A`qK,g���8(�6�q� 7&��F�z�+��M��)tb�|q�9����~�����T?F�ɶ�~9�{q�Y������aq�[�3��]{9�lb��&�X�Ҳ���8��^L,���	I�<j��GM��g�/�|�V|x\��v����e&�N�J���%#��}f���u6��6}�6#`�M^^���mq�S��):���kB!(eoIZ�H��i����y���<�6:��QL�,I8�̳�Xw��:a>2���'8����i�ok�+��]���G�x7@�=�_=<!��%vG����+O��ӈ�Xs�yd]�s�`���ą��XS�gh�(H6���-e-7iದQ(�H���!���fD�A��b���G�l`�M�/Z�_` ����1Z�N��l��t �]�5` �$%�|<���ړ����{>�-�aQ�a��Ő��Gs�M#�<jT�rcvX�M8�H
ń�Y:9Z�����*IM�=�(�g��󗜼�}�ϑ]B��G�ˬ��M��e��Iz._FA��A/>�Isc6(Y]�/�m��X���� J��d���j�LjS1�H,��*�aC��ּ/��o���F��E����c�m5�!J(�+D6��ߎ}Z+&2�V���e冑�	����2���L1�9y�3=�Dy�k@I�ӝ+�Y�*���@�S.�D�"���u�2"<^����
xėPl�el»vpz�+5\O5�[c���T�6)�/���GX�%������ϳ@��pĽл�6��_�cpe�4��_�Se�jܾ�	���5�} ,"Eڞ�p��&����~�ÎR�Uaï#g:6��g㔅�Ǹ����y�^X.� ���iY}*n���"#JGT��)���(>��gV/x��ǟ� U)���Tqdhm�k���#_r�x]F�%Mw�������Q����"�ўȽ � ���HuҌ�ڐ__���n���)��\h҂�ۡȖ	��g`���n0*ӌC��u����p&�-1g��e�r��o�]���7�����5|�F*��ԋ`�'z��-{�|�8<�&����3I}R?�v+ɱ��%�!�3JQ�u#,Zj��84�(��f� }3���\{ 9<:ՋD
��0^� �G;��Hb��?��5z�$R!XE�=�cӶ��Vlc���k���M,�3�+�Ekzd��k�_l�(it<E�]�P}�
Vg������ЙˌC�F�]e�U=���彩�f�W'�$tt.��~�"w�̢��s~\rcefX�uzwS�:j#؉�nt�E6�D��=�<��i�Z�0D'����B�w���u4��v<VL�o/���"����q��_5n;E���z�/�?y���B���3��K�pX9�M��H,X�������\ ZԄ���П�򊲚=>��+���"��iW�q"���;�׸�p͋&x`&�28R*�c�c�ٓ=q�7l��YD��tZZ�b5�$RG�\���z⼲���s���]6n�2�Ӹ�gɱ����*C���7�+��`�#Y���-���eN��G���p�1F=cx�2�}�k��69;��G�Sg��ٓ�S�T�f���ķIh�P�2 j����ٵ֎*�ŗ���!.`��ψ���x�Q���T�5|F��֯u��nf��E�0dW/P4
�}ȿM
���m�G�*N @7W���ȱ��5�!c�8*��x���\�4��F�'v����"��(;*�>��s��5�K�5��#����e��<���{������;��@w	E��r>@+t�ϼ�0׉Nр�7/c�fܘ����J��p�B��k֥�����F��f�(��x�0"�^A�֛� �Vi�%�xz=jr�	�jG���?�Z/��qh}�x�ufy�Z]Xr꭪2.��k���zԫ�_o�/�+?o�4�feϹwPQ�L��K��wi���[��)m�K��=��V��5�����Q�)k{_�Q]�z�s²0�Y����LߦUo2�6s� pMJy���Ѯx���h�Ņ��	jF��?�>���u��^�,��~W8�
�� #$'"�g.F�x_��	ǥ��e ?����t֜���b�� n�gT�[M����߮6p��v���ƶ�9
<t8'��̩��}��\%��z[�j�{(����5I��λ�uT`珷j���\ݿ�F�P1y��Z:�ԭ�����1w���>$���z����_�����I��M���-�-��&�wZP����÷&C�u��9z ���O�b���9��>?a�tF=u�t��Q�h�C�E�y�Ժ������%���A���,i��mF�y&�ND��]� u+�vy$T쮂�q���K@��1����>HOS���Mуe)럌�<p����u�ǥ��		j\���8���̮�oYt��!�(J����;h��]��Q�X�|��
��Gm�zn�aF6Ժy`.�H�eM��)p�`�.���П�~H(B,HBf*���n��p�����wt�К�۹��}��C��8���M�t#���t�s��Q����D
lvF���[�f��=b���g$ZY��fAК�[f�8H�"D�^=�BJwh���ϻ�p[�4+�0�ʡZ?e���̩ml��K���C�ZL���e}����w_y,mI��q���5)��D��<\�uG��ZJj�;|�5���q���Ieu���{.�˂����0�n�A.�H�dw�]\�]�}aP~�ǧ7�������+NH�Tb#(R�����Cq��7�+3��g0���Ë���p�lA ��:h��b�OPz� �;�f������Y��۝���ῪM&P�ɰ��q��:�x��'"e��e��*ؿ U���`]��JI$� УDzg9<	s^,�����TL���_#6*�B)gV�%�ӒTe�5��G�}���_t�m}�E�{������o�E���<Bu�����}}D�0�x���Nq�M7�22�����^θ�EM��Q�oG�)��H���i@��=f�ŃZ4�:<͍g8ס�SO��6#�3�g���|CE���E%��8�ŗQk��/�&O*�9���q�~���[l�r/�}!�m�BLig�n6o����\������U�����`w��y�2	96~�D�J��_X*$%���>.'�󍨨A�I��F��o�5U<֎�b�Kb��`�e�/ĹjF�e9�F�"
�;׶ߡeF�G��#�˩&W�Is�%�q M?$Z3oQ[_�_�;qV��cp#&�ba�h�"y�b���#�VEu�u����#��\�w��if8|�ȅV��8O�z�Sz�V���qA�7J�]t��m�zx ����j��-�eHt횘[p\�2��7�k!{EQ+t6#� �Eq_K��S�D���J�A�߭ �3��H�`���j��3�Ǔqu�7�.�^��&����M�]���8*	]�Ol�p�10j�#���}���8!����qL�[�kȬ�쑎��5Z}���EcJ�.�cB% *���,�ȵer�`�0fk����$'�@�����-���W��H��W�I�ۡ�b���e�x�@��aM؀ǧx�f��I�^'i���Js��%$����_.y�~�!<Ƅ�ԯ��	�v��f'��d��l���H�-�*�>����}���
�_��ECCp��e�&\�I���?���0�9d`c�TڣI$�ާ��	
.�����.RE�I�`��ML��q�P^�.��/켕BohK����+Ios���E�^F�p�������	8��B�7�{�����/���1�^.s
1B%���Db������g4A�Ҿq	���,F��z��0-m���qPJ-�#-��ut9�T��?UM�kt��X	 �%����݅,睊��I���/���^;�7�dU���_�� ���U�i��ȗ�ޓD�'#;�:�I��>{ �����9�k�Z���i�.���N�v9ʍ�.�4��1Ԟ���p{�m���_�t|�K�swm� ��;<"9�R�n??1��d"�a���.=}oj�Z7���5��$$���?~���ay'F��	� ����)٬���bo��I|�^R�@x�x�(Xs��QC�͚�C�u���T�Fu2[�n�B!�Ôh��hru�pi�JW5�0��\���K�,��2����7����<`^��G��qÌz4�8�{�-�00��E[g�	�g�-��d��^va����ռ�&u3�	�,�'9��Ry�{
�<ڗkp���ۭ2L�(��2Qt�7��Sb��("���G��al����N��>�e� �Zj�����Nk.��a!`t^��}sd���ۯ�5��t6����{Ĝ��y�
,$-;�H�Q���,���&w�A�O8O�K��@asܳR���D��h~�NV�K��55��w�Q��'l=c�d��T�:	�W�"Q[�C7�F\S1���xN�����^{[$O+.�.{�Q���؅s�ɯzJ9 ��Ed	�i���O�As�s4�#�C�)Ia'Bx�|r�����6���D��I*,��o�S��K�c�`{�ϙ���d��M`�"᠐93o����q�<��K�AWA�)LM�7>�N��k_u�N���S�Y9aԃ�5� �R�o�h[�V��<�i�#f��	��g:��a���.յ�f.x�!� ���X:� y@�W0�U]O��g��~@�Y������;�A�hj$t�a՝I��]]iV���J�rE�0 v8��VF���W$U���-v�L���+��}9�S��蟮�BV�v�� ~"�}���:F��z��J�!M6AI�dT��z������x�l&�3�^�~����o��9e����:"�"[ ܯP�*t��ˡ�+d�p�mZX��^!��SI�����=�Wh�g0�tъ���Yh è릷�f����������� ��S��xP�U:ݨ5�>(N�'��K�X�a�O��
�BEn$��ҝ�;Uw��ؚd1ՙdž�5��)Y��ֺ�7 R#����{���ȣ%X�h~��=��x�a����*���j��jW��L�vf�������)��T��r����E�V}�!m4@t�ʜ�8P_�9�ݥP��͘�y�#b�������P�q'\c���i[	>���Q^X�J*S��d�J?��|��84����'�oFf^�m��K�H茄�k��9-��?��Pr7r���V'�%�}mCR�:�F�F&'�j_�n~�>"�v$�:��4�%��R0�5>�%yrJ�}�%&}���ʅ���s����s*ꨚͦu�ɥ;�,3�T]���6�Oo�v9��������/ �l�7�<q�ছ�wR�Ұg��	M�����Qj��9���&n/��˕�%�=��NfV��A��7gdW��G������[�F���p�=�\Qt����F�*<r��e�̜=Ή����2n�E��m��^,]rz����v�u����u���U��mI���{����RxVl�l<z�B]k)�6�خ68C~c�cqk-k��J6��S����s!
6}��J�ɶ2��s�f�=Nb$	�nBpU�2O]؂���˔���s:�̯�P>X��h��NV�9�v��x���':ۺ��,��3�#&��q_z��*� =ԩr��+!��eB5�"�2���H��^�b�N�,�l+K^n� g�
HU#�9�@�k_J�\˿��g`7�X��:����`�x��[�ntb뻊��nÖ0�+!��h�l��&�N�x��4�R`]�~��㵘vTv@S�����o~o[�����},a�7�`����Yp	Jp��?0�(����O�ô<s����ED�����I���w���AEji"q"�;�E�D����a+&�8��DsB��f��Ѳ����3��S_��1��!CTjJ��9�ؘitJ�J'�S��2W�Ә�m��/��W�@	˸�O��Ed]H,*k�֌�<�W\]����s%����g>ap���^2����`�����g��:���7����JH.E+��9��@O��<��f̊]���O����ga(˱�I�f�A���mrg�f�NdS��(�mX�Ά�	3��7����A�X$JL(�������c��@4�ZHX��!�i����b��:9�.��Mz���0���9��{��@�����Z�s ��uR8�F�6B����l2���M*���wxx@���Τ�n�%܌��,�m��H0�"�*[�M�����"擜�~�ϛx�{W �3���	Kf �[b
lXLG�V��aR/��5���E�ƾj�Aϟ��I�E��0x��F�_��F����v��d(��*%���#VbEq�j�}�fS������1�!��zO!s+ŋ��*��X�t\6��D�r�R󜘷���i�cL��z�
���}B�"���*{�P��7I��t�)r�O)}��R�h��t�Aۉ#`M�j�o]�m� ��ZU��S=��o���k-�戊��5��,��H���[�DZ��{�����B
�ƜˍH��RW+@
�g���A#��]�9��c��_A�����rD�#F�L2: BڒB��X��p�!�Zz�K�*9�c(���Նp�pR�����{(�b�&����W�i쵽�w=�dlG����7����_[�t���vU�|b�5^*��T�,�9i�����X��v*��i튔a��}�*�\���ƅ F�+ �{�,�Gt���V��E�Fh=��7��vi��h���̓�N�|Km^(jՎ|�v)�n�_�u�Q�N���D�l�o��(l��%~`�]�Y�memR��VnW�?vl��`6r\ D"�,}j��rpE�h5^�h)r%hz�i�f*vAgy��d)t<�L�Yrp�l� �,���b��A��͚�$ ��E�"�(E'�óG�a2�J�hZG�λr�@`��p�N�u���s���]w%.�0�Gh���8��r7EȊ7��nl䜪d����b��Z�HD����3o�Qd�A���U%�ap��z�s������|SK�1Z���)���J	'�4�B�n4m	���Ƹf��N3��v�%���]���]ގ�����s�Q����a�.��w�����y�.D9�Hٸ�5�8$���,n�I4m�S���G�;�/� �Ce��- p����������%�a�W�2{	��+P�k����g�nf^Йq_��&[��aO�N_����R����9:�T~���.A���O�B�IJ�=5�C��\Ø��P_�A!�:�������v�+P}OaOj��5T
�}l��Ї[N��b���/L��'�WT�0�P���|��M��sD�e噙�汑lv��t�Sm��S�<g����J܇�22��N�'"��W��P���p�n�[�noAE�{�y ���aˋ�o5�CI�^��'��&�����;�TX���q�6���=d��'��9a�{"#	��n�����:�w�H��X��x��y�q:���'��{!�Ա$וȂu���#�`p�Q���ӅN������7	S�l{Hc��n���2��nE��Xp:Nko��+�P�h����R])�H!x�{��&��̩�����t��}�0y*�xWyΧ�c�r�=hXa)�*e���H)�1�;�g�T>ځ ��f� �{��{�,z���M��Q5�\	.�������+�Mޞ�:�AA�HH��`v��]ׅ���y��/�Ҙ��v� ����y!�:n�-��.��gҔ�(/\a"W�¢����4��$�)H����!t.2M����/P��F@���y�g��ԢZ}�7���
�W3�fx��~x��bJn�̛'�� �6�����
@uB�M�mi�A�)���W^k�����.��u��ʯM<��uK����3(�32I_\�	g+��QUȈ�\�Jw6v�Z[��eF����+�]<}���[x6HM؜Σ��c=�l7��9\��O��73`�,��"�su�]w�*�/_-�F��x����&��]�Q(v�_g��K"|���9���0�M��s�w�2(:)�ћbz���� �Ե=q�<);���ا:���ħ�[2���JG�*��*���ʿ���Ʊ��&t���e�伉�s��xv��৘��ȋ�tP���^s�c|��|2��P4�O[���am%���/��]�g�y���Bġ)���y��õW�;Ǖ���˥��*7O,t�Nݟ�%��A��2�*D�<5Is��Wu]���z�Ι;����U�F�������}9�5ؖ�Ը�	�#�,��Q��&V��u��F���H�Ċn���d���I��'ܰ� W8N���FI�Say@�����t�D7�K�$C�>n��~Z��(�/��IV�m������Eb��p����W�t1g��kf�w  lM�?z:�.� �*k��e����N��P:���RN���4Ed��T�he3 �J�����$�=�sҎ��_��y��tNS3ٽ��u�SW��M��k�QQ!�m�X�im�W�ݦ�":sd>g��T�̥���M��p#C��8���4��%�}*�1޼j�
�k���J'��ן��d��C�Gu����逸�'�����2?��	ߋ�ݐ�j�pΗ��&�O��j.��;cJ�`Ĺ}��L���j<�qhX��O��J	�3Ќ�$$/�|�����(�M��^ �t>��/tp���)Y��-��+1<4?'#5.�}��T�"��)�b�A�
Պ|`�nN$5>���Mo�eAΚT��Kˡ8�������X+D��8��
B��P��Wl�#�"6�x#��e�܏��u��G�����/_��<���O@�PZ����zV�+��^o�S��~.�įƫʧ6��l��:�N�h�u�w^D��J^�-h �6��/@4������%nH9@�~IHf�TDe�B�UhLv@��K���6��)hH�gcK�#�T��<�B��t�u痧ǈ����#�� ��Y�98�Fi}aBH�a�^�kr��S�Q��uϰXu��C<�3��b??����]G⻄!�6�b���h�;����jr�AP���d�|̾�t�3a�.-�����%�UBwjv�����7�qS��5�����T���w�+a.�*��9$uÔД\� ��>�0ъ;�
�Nn.�h��L.ȭI�ej�$C���e`.��L7z��&CK��T��$y����ؤ��}�X7����a��T`yp��e�&Gp��smǀ��|;����5s��]�c\�0���m���fxg�������<hOw^��P��>G�#�ɡ %�OJ�ek4V���,����u���$��5Mm1o�?#�!쎍�j��JP/��N"�oDQ(F�>��Ì�i_�� ._�P��Ζ}(���Wڥi����͙�^���N[����e���k���D,T��)FN̎��AB<|%�N��~�F�b Mr��w'�1d !�>�GN������<2(~,�Sr$�ry�v���G	ҹ
�&���o�L�:���q�3�	:��5���A(5�q ��E�'���]�jPDJ:G�q`hcSBT�oj5e<e�⚘��CA���銂"vg�Fm� �%`f���y� P��� �bM���u����3��q�{�|�X}/�㨠��	�W@?3A⹍�2ucWƱ���'�[����'u�sa�2P�jva|�F�aJm~��nOцBc<� �,��"�X������mo���C&�۝��=�nS�Q-_���m�Z���:`ru������)!��-ꦩ]�`Da��!��Y���Ω��᧟fW�X�OuWeUe��ma�L�JDc�Y"�$|���騽+��]���d�F6G�#=��\����U��&��h�T���G�y�����ܰ��Ɔv��@���Wi.�	ؒ����=tj���)3��ܨuC�}��I5Dt���nB�qF�$)7c��6��8���ziˇ1Xا��j5.� dY9�2�K�Š,A�)9+���0	����j�1Lr]��oPx����-�x�J~?m�h�L\���o�+��vv֌��s�w,�u����W�bU�B����(z��b��7I&wa�E��)�m�"1��E� �D���G�&�E�-�$
凥�[���#����@�BzN��N�xF�A��\8�>m����c:�GT�ci
�R*�y`��Y��f���y~�C�5�InXZ��;aZc�����<f0�i\�õ̐�x��Z��j0Br��&w$&,�ˍ=����A���DH�+om��.,H���[���H����O/k28�*�"4�n_%��)bvUۅu]R�B�=Ano_�ߊ,ʔ��E��O����~՜9V���jh�?]����(��=��Z�W� y?���mO{���������s����`Uʤt}:��)�n���
�@�	t\,�{ĵ�R��+�{�Ta2fIq�����f�th{�Y8�/ȷ�r�x����}Z�JzD�o�PlS�Sy�mHOO��P��ecC���뢞�Pk�},aѮ2�Y�5g��h�J�xD^[>^�Q���OsC.��F\�%ٽ��_�^Mj������cd5P~+MC�-U8S�
��B2I�ց���6�zk=G@z�������f^��@\&+JE���)�=���`&jad\� {P�j��EwO7��҄jU���/�$PO��]�BZ�Q��L�i{��aR\�?cs�J����J�N�1��#he$�-	�ֱ�m��\Q����D�`�S�"�	t�<~�鮮kȤ��|o��g��P�$~ݠ��|����i�S����cb-�m5�y���I���E�l{�!� D�E72E�S�-��*�)���<
�C��J��Yg����L�,�"��o�������Wv �@��@4uM��WZ�Y7�67-`���*yq0^�_;�eRмSX����If��P�9��Vo�T�Q�>�s�ZN�X��{Lc��@�N����[<��MsW����M�C�S�o��N���c2����h�����/}��)E�ȥ�UQ���,�Z��}[��*` Xڮ�#o����5jޓ��*L�����q0�Y��UX�H�����{p�,�؝n_��}�����-������Fϲ����������\��F��>���fr�[ƅ8w��KG[�}YqY���D��a:NP�ŠȮ��M�_���wO���c�|J��œ�qw���͚l8{q����_%�c�"
f�-w*���ё�<:=W�WHVΐ[�f�w���x`�Ϡg�VPD��o(�)�.uy+�3�P4�ؤ�
��0Tì�s�D��9��u�����	�>`�F#�§4櫉V��iC�va"�F��ĈT�uB�D��9J'�Lkr��+ �=�����\5�|��x5��݅�W[%}��PJX����D�yl�b���t�HB��um�ӧpPj�����=ƪ6��O)���D`�I�zz7f�`��=xӽe+Α��囖�bVS����f��ڼ˴��:k74V6�5�/`'G��kB@oX� 6���)���wx����L��u��}}Z�g��h�W����[�����y�ȳ0�K������g���A��;I��Dz���G����C������¬��~�w�i/�˭�v�oʇHэ{�u�HDYȻm����C�ʍV��!�{k�V�m�]H{
/�o�T_%�CeK�����*���F��a���V�3ݚc��7���i��{��H�~���+�H�(=4Qa������r��w�Փ(�[��	���h�k�|� R���$S���ܥ��/���d��j��q��̭�h'����w�YP�L�@��/�&
�v���ÒZϰoR(� %�R�6�[^b	[i��G/5 ���O�Vl�A7����<�8$�W�����`
���*���y�����������Z�9�Ek����P>U�
�������x�o�]6���3�������q��'����4��'�����+�嚂a�<�a�*{��9����ާH�I��y�k�7f�"��ߚ� �����N�F�"p߯~��	�B"���7����Ժ��.�'<�j���d40���������/#+ ,9ֿ�Afp�y1�ի>@�������5��V���`�f!�ޖ%��AN��*��r�Rd� �q	(��R�Q�`��Z+���B�<�e�o����¿���6��v��d�r�O���%��=P�J��nD�=J?<��i�@��]���.pYE��R�.�bR�}\�B�,�AN�]�]��M)8��������af$ZAH�s�Oc
�j"��)nZf+����� ����b7��&?��Gz��/��e3��s��q}�1�0�8�<��d'�|�r8�S�����q�<=+}^���-��v�vk��O=4[-�NxL-��PKjS�\G-�H]�#�|�qZ�4GS'Ẅ�^�}�����`C�qXBJ�G�<��7.�u _�Ȍ��P��'&=k���^��.�u9J@!��C��p��8�H�Cb�S�I�|�@BZ7�aT��-�[ɝr���;V��
J���o�g���F�����v̱�C�i�e���O'���?�W�����_�����m)m$"��n�	m��4gb��Ȼ�}d`�T�V+��#��Gw1E�x�6���c	��@,3.��<{R��nU�60���Ye�r�H�{kݨ����.�G���fV�A����)��~M�K��-n"�9�� *:��AQ�}SE�p�VՈE`�o@���wv �����^���Q~|T�k�:�LA��?����y�M#��i�J<'�!HZ���_�݄�K_�ݿ\8��a5���h֪��p�Ơs�&?��R�_d�����N�=��㤣�������:¹�� ���fO݃(c�6�{Ud�<�X��EA}��Ȳ�h�{:�@q���֤A�6�>y�x߁;R�r�|�@OMb���o���f�2�p*�����00�$�bv窭���6,�R�Tӟ��rɚ#��H��_
a���ͯ���F�f.B ��B~�X�l]ll�<�������A���\�ˌ�$�x!)�yH�){��o��N�o��^ԡ�'>P�>0)ug�ۉH��\�ɛ�/��?+�*��R�[�F������%/�7?́}Ѡ��c��Ø��$�1��T��?x�TY���W�I� 9����\�&��x	/�����'&�B����Lm�$-�}c��g9�gy{ޥn�3�db�\�c����#�8gJ���FT/d*R�m���`�f;Gᴺ��Y�J8�f�p����~Fg�Pr��$�-=�ts���Iۄ��#&Xv��S����Vȣ��`�VP��w�����8�!���d�� �1�T�p�q����4���l �3܊yff��RF7$�D�&�O0�kF&�"T�^��E}NM�]��Ng�U��)pf��B/���
�Bh1��>{��n1"X
�xi.�3"+H@	X������+s��O
��(�_A�����X�>��{�E�LC��jT�?��YU���,x6��Fʾç1�#)�;y��&�� �W:�E�{a W�G#Rx�p,�z�|�a"{�p\��m�2o��ڜ)�zE#iN�i9��j�o�@�:=&�>(��8O�n?���i!��)��Z��5Ts�ŏ��H`�EA�ދߤ�d�bW���T9�)�J��i��[�k�8�7�j2?�GX;�fi�fF&�mT����I����XYȝ���p�mǨTzh
���k��U(Kwe�P���S��h���I��3?�#�I4�C�b���6�砫Ę����Hʬ�MMzE�����
U���ݕ�)O��h �p��HH���cZ�0%�_�G����4�R�C�0lf���D��j���`�e~�˯��b7QN��|TH�$��hSj�z3������k��?V���&�25�e�
��u��]�h(��%?���^��	�Y�ڸ[��UWY�3l1���@�5�4��+mo�y��F;��J��?�֗*#;f��x�q�Y���6A@E��u�q,�{I�b��a��N�Zvڦ��-��Y����F=���]�[E��*`�:��ٿ���ܝқ�u�䁩�!�9i�TA��� ��.���=R>�r��K��̎��V�Ra� ��9��e�����r��sp�ދY��H���%���L�3����se]�	MF�y�`�����G?/��\�9�,��{�, �h�n�,xU���]�zN��ˢ��Ktn�ɶ�����s���|D���q��㷛��uf��M�~q'���8wg?��'�u,��7���C'^+�c�<�`���\�hK_�L�"
�GU�z⸰Kr��n��L�7A�)����U�=�1ˁ:�Ec�����
��(����#���Wc�������1ޚ)�I
�/��\Q��r�H�iO����m|��z��ZC@�@�a����$no�h�*'���?rB۔�nR��jK��]�~���� Ҫ&��i�RL���7�V ��`%�y�5�Fih���j1�,1�avҒ?I�l�^5@����̀�_/�NO�yg30��f�=~�˦�Tu��O	��gG����k�:(4���/��_ә�L���X�̴BY+�](;����Z[ӣ��ui���	�8"#
�Jq{�.M�*��-�پA�3�J��$�ZP��8�5��^Ut���_*�e�-?/_�K�h	�.]-�ƨ��AƇ9���ug"���ew� /j��I��&���;7��a���θ�M2�ǜз�����RBx��������q��c3�FBL�&����B�h�pI��?V�����O#~�j�'�{��Pێ�|��7���� y[y8�����hA ڞ�|�R�aGn,�p��k��� ]�P��>@MU�129$��Pn �V�G�?O�����V��;S�fW!����oD&�� iҚ,t+��8�2J���W�c��$L��1Ya�_�yJ�����?�+7%���Y�l枆q�I�tc�]���"萂�JyGk�*��~�"V[h9��5l�˼ķ���.��i����\����V��h,��w���-������V��=���ߨ���-�j_8��p�+.�=�3燸����h��@�K�jn�/���1M~�Jan����I`M'�?sZ`�Г�n�5X��X7{�g?5�x�^�c-�����O<羻�Y�V�'�����̝�U�^-Nrz��y�ͅp�Q���ê��4����sx�Jk���*�}/��{�bjo��(0L�fq�c�����K؏��HIl-�t��)w�"������dL:p��^QS�ۇ��݉��J�6E7b9��e�,5��[�eԡͥ�j�}-{���>tǊ���Ɂ�P�~g$���^B �p��JڜJOjw���;������Q��һ����@�h2P�sׯ�+�2{/�(c�f�޴ѫ|D��ѽ��?װ���w��[PN�Ϲ�؞&��b��\gp��S̾�$,:!,��b81#3A�aN�v��2)=��T*5�ZA���E�F��� �D~���
��g�
�q��#���-p���6%��
*�qJȂ�[2t�1�H?`d�>5��ek�԰�,��Y/������4��G��t��C���Z'�G3���M�LsrD��R����3��Kls��3�A3�o�P�&�����i�j��i���V�3��Z�ҵ�0����2#�[W��2Xo�K�+4Vj�bd6)�� +��%��_������RϿ:.���ST�ĭřCR�\�M�ᯠ��K��+O�f�M��0�C�)El���GA�x���PF���+SZ��1y4�DA4 &T��禤�Ec��k�q���K�AIB���.6�4I�5��!.��*Jd0 �,�ç�Lo��IԙG6�z�`'�_��[�	�6���WHt+�?`��t�X9\r�8Y� ��s1��c�����.rr��m�ɉ7������`�����"Th���ҷ��&�N)-L��ޮ��J6�="��uG['nG8�e����|!X�;B�z�$�(*�����G�Q��<�"���|�����F��ă���w�~�\�_�w�:6��	�ב�d8�LV��	B���a�5��D��=�\)���)I�C`Ю-|6��w�R~d_;�=��jc]�:�����İ[����u��5�.[�|*���մ�;�Ebо3�����r�.�U�A#�){�(T�?"6���-�ӿ����".�;��g�As!D��k�� ;�N�f���c�C�
�SL3�y�Bp����E�w��ģڐ���v~��9���i8]���%�(��z
&L���{�oƤb�e^\Zx����V�iA��r�6Tt�%GZ]�(��c&@a�YI'��޸g6�L�f�寖X�R/��4����i�����yD�4O�`����zԀkɓ����uX��U��|	���$HO���]��'�{����Q6a�@}F��<�h�p! �卮� �?�����@Up�JG-����b>A���{g���;��%,՝ut$���h�̤�
{s�`����������r�ϐv�W.\3�`V��7�c��M� k�z�lHp���u�6�dt�00W[BK����}� @�+P�����[��Oc��ZF��������Q�1�p�Ivts �U$P�Iѳ��=��73��2(}�����.TF�ǃ�	�^�]�X�W�"�[s�����o�D�Ym�8#�/�]+-kNU��
$�f�D �m-�&2��D��/�z��S��@JO�
k�-�q�bZ��L��14¦����$&I�F������u��6 ��*^=r�0���^��6TC;�G��:*�l#?[��L�&�������:����]>{s�[�oɨ���@���rq䫧)���l���3O��}���~�dr.6r����-���Ⱦ
��|T���/��\�r�4���mFl��� ��ɏ&Z�.ʃ���?cI��	
��ɞP9>ڌ�K��i�?��#�WAܝVW�eR~M��T��iN�I��>������UF\�iW��I�&�[���+���X�������%��b��]"I���ybՓ��h4�^�V{�[��ֺ$ō��,�b��8�C�*~|�E�U�����Y�a uL/����tpjx����)׈x���Qx�ƹGV�?:F�Iz\�X�V��y-yESw	�Ѹ���gP��<�u��Y��_+^&Db�(o�������n�]�����`Ws��<[r�\D�lW~����Hp��k)jwc�n�D��2{�djұ6����/�����}�"@�N�;-Oi�$>���_�2QBÂ]��8��{>^j:kSrH�!f��E)��ѩ�nQ0���N�@e8ݛ&p��/�mV`wJ��7z�6�$��I(|ɞg��^>����.�ѻb��'�e��M���?o��p\+@�Ц�?�;��);��*�������P�8z��:Jn�g�����y:Q-)8@����S�G�ݬ�
0O})7a5Up�Qe�cu�_a5 |���'�4�4_��J�z�=��uO�0��O���U����Q$]?hq�M�m��Jg�1��,�V���\NX"V�)���-����S�a��L��j5�4�	>꜍R��}Le���c�i�Yþ�!R�l�F�oI��V��	��@@f�%��sFjǮw&�0�&�gj%"1��"eK83�[LYw�����/�!Y���uY�"�`%BlD�����M8 Ѓ�j5l!�W�AA+�q�ܰ�B9��_'P����ϾS���.پb��x���+]��>:�f�~�%?�Pp=����wm����]����QT�*ݱn|P�V'���ې/M���+V��@��᪠Xq�u�_,XVPr����p3>�<D�"KJ��R�	����[콐k��F#���T��E��W��1����:�絙�v�ZȎ>��\@Z���$��ϡm��H߼����\� �`q�]�u%P��?��Ad&MlM�\��0Oo�X�'\�]�I8�Y�����".�p
���G�[���Xf#�x��O�D6t����>[������|8����I{}w��1#����6���QD�$�����*������G>5dg}ڸE���`�a]�jD���*^M4��aa���V�O/1ƃ+z{��涫�H7v������K�$�2�*-}�����-�r�����#*R}w�ɏ�e��󳉅/�C���%߬m��ߦ1��n��Y���3��)�R��w+5(��f�t���>�Ԅ���[^+�C���2^M㑗|�u'�~�<�R�\=�����g����DGE��-%�t�ꇐV�󂽓�ݼr�`�Rt�!Ȍ ifӑ��y�s�+d�Q�*��C�?���]�u^���!���$~/��@q*�:�
�7&��W�Q?%p�ȇ��e+PhH�U��! .+O�uPa�Y�%���7�V�I�SԔ�]:���X�5��,������_�*��6��zl����MO�Ge�=��{��!�DI'ĥ����[�"̛'<�oX�c�������{/�A(�s/�BC2x��ɷ&�y���?�_���0b���$��+-�,RO�j}�� ���5{���W!`��`��jRĒqƷ�2����!�Wm����$m����(�*@�L�PL��� �kO�Jy�c�l�K\M���=U�6���Cl��eoL��v0���j8�L��5�P"�v��à%�;�I�0����YF�l����c��l
q�}Z��
��A�M�蜸��ݱD��N�]I^�*� ����z$ K�9C�&����=E��0|��o����
���`�}�]
S��>a�~:	���yK�3$il�{�`T��9!��kbk�-������G�oēg���(��s�z��$_���喵1�����%,Z<=,�ğa!'��d�:A�r:���#Hdb�I����~Zm3쎬7�8��Yv:ʎ��M���@PB�=�Ȕ+QgM�Z�c�2�:s���y�|̘���lzd鬁�~)�z^V0�ϛ���f�5�]��y�m-�WIX%�h�I{�^@���m��6m{&�xZ�W�)*���jA��{�B���_�NI��u|$����]x��޴S	�{A^����蘌�ȃXվ@��v�o�W_��Ee����ȇW=U݇�*+��x��	".�:��aE�V4�D?�c�G?�J�L�#/�X6ܮ�Qvkc?�Y��$���wk�w�������W��hP��B�`w#:�bYM������i�(1�I����6�����/3Y�Q������;a��5 �+�ӿy�|�H��}2]8�'�����C��u����Ǹڀ�1�#�Ƭ��7�0�1璏!������^@ ������2�[Gd�M_��pO�	4xʥ=�^�cc!	N�\�a�T�lF�9��¸�t�c�D#f,��<�i|bS�:�O�վ�؀/r.x�Xs����+.�A�e�?�vK�CoZ�'2 ���``[���A�yt����b�T�h��\��)��=>��}�gz��[�$?���<�-ԕN�LA�uTL����޻����K�Bȝ<Hz>!25��ޒ�θ4<+7{���iT�+h�I;9GpyO!��ə��]a7�����L�����,���Q���Cl��B+��i=f'���X/Ώ͕U�*��v����%K��0�F�a�k�\�fnWR�+�A�x����W�f�@�N�*_�eW�,l�,�Y�[+��� �xI��I~
�Y���`ے�g�8Ux��.5�R��*i�O�R��s�z��(�7�����,�<�
�+�Z�x�o�%���� i�p��=H��������Dp�@Ɗ���ux&�d��өD�u�P�r�=|Cp��z�6T�L]0���4L)�ʷQ ��i�S���>���*���b0-.�)��4tdE{��X`�����Ɔ�B^;�$P0�@;$s�w��o�{[��R�93)�ʘh�����췕���o�#:r�/���y��û�J��FZi�n����+�e�)p�É��7)�PSEP��]m9T0&�K'x�
�8d���Z�������f�P�q��A���u�+�� �p����uǾ�����pL,n#�r@��a���w��vIJC�?��4|���?]�I��m+ކ�ޫ���ag��[P��� =��� {0��/�+�z�&2Dx�����n��)�0��\�]|��_�h]�����<��9��~N��;��L��H�*f��?�	4yۡg�t\M��G��J�
�V��Ä�����"� A��bk<r\�Т�I��^E�:G���w�X`/������G�gQav�K��J;r��J`��l@�@cV�=�Pdc�Y�^>Yۘ���~������:�
�����Ie����
H��x�xˁ�e�*B�\/����v/2F�d�
=�t�F�,-%�3N�rK�o��� 3^P�ߛ�p�FX�����)7'�S^x�e���,��D�|��@RV݄l��F���R)��C��]�c��L�Kf��ko�D2v�EY�S����y�\��!}���	겵�#XJdŠн��ب��8=ԝ��q���X3�3vpK���g�Z]����='�:N�dB�j�>�{�������K�Z�oF�$�֓�"Dmg&S����'�[��ⲃ�v�8�R�k�i�y�����~ʊ\MHQa*�z�~���E����aa�Y+ds?=��k�EJ�ZS���i�?�x}��_�sχ5���C�VE�^�;��Z[��ژ�l��ƴ�U�Z�O �ꃣ��wL��N��B�m�	--�AɾhKgBnŖ� )@*�b�8NOEݾ�e9��#�|��H��;|�H�B� Y�i�9�#0��q5ܗ�Y
|	CC��7��Ա�ˡs��w����FDL�d��Z���h�sK�=�;?L��`x�ú����/�_=�)z�r��>ò��+�E����`4���e�*`R����f�� �Mڤx�_c�h���L��r�� �8�	'�eZQ�~a����I�����~��l��'E���xo׆��Y����1V�N�)�<$����f���H�f���e��%���X�ݡ�d0-g�
�8O��B��
�=����M�g����}.b(�#��@�AjCQ\<򪾐S�QϾ^���˞��3x�j�}y��on�ɪ����j�ڱ�E���J�g�$]�!4��u�ωF���FA�ݖv���P2�0���S'S�A3���PZx��n�X� ������E&�t���M��7}2���%s�K����'Φ��?�t�Y����rk�X7��$������Vֱ��?�[�ђ����#�+�����>N�(��ve��i|���3�3��=ە=G|»��,J�v��8c��ls��E.�Xvm�Y|]�l�2�� ���=ݩ0��zf[�S+�"^ڍ��ôb�d7��b�K��Ě<D+�2�r08�����;_�{OA_{J����`K�D��R�M�Cc�|���Si.awP:�E�@N�%����� ����鋫�S��4r19��y�@Gq�:�f�{�~L����ZV:�C|)�7Q�D��V��9	��}���T��S���Y1����v���	�,D��Ѽi�.��O��X�>I�G�L��^\E�(��t�oT%��s흆����g����� ��ޠ����$YI��Ts޼��g�iU��ul@�(��dB�����Ts�H�[��~�32��5x���H$X���8r1Ø�=�|�R�.Eэ�5��Z�"K`
���1UWf��zz m$�� Jd��<ǧ�7��L�M���@.�7������Bڲ]ln���^��wL�~��ͯ @m��CX���G-Q��d��/P��л?��.��z;{ko	�jĞ��oOSղ�"v�p��]�p��� ��:�����{{
&�٣���!��[N�K�sJ̔\�3�;¤���34Lt�N@���߻f�,N��h?_I���5�}���^�z/�m�>�+�͑�RQ`�b-��IXr��HS�
��ߡ��꬧0�թt��`����n ��T����=��7��vi\�Yv`�R���[�,F�J��̽���O�� ��v��:%�J`)@yC!��mu���|_�I5�������Hk�t̻l�����q�9A���;41��7&��`��bi�+�� [6[h��/k��4}��SݒJ�л5ܿC���=��]�o���u"�;�F��n�0Z��m�4��Cֵ��?�s
�:�4��(ݰ���S���XL���Kw�B���~�rEM7@�P��/��}���N��>�者C�:ёɆ�]� �k׉��c��!8��A�#\ �"b��2/��nm��O�An�6iz�Sveo�Q�e�A�6���CI�#���wc�JC�4�
�mh�>z7:��\[g��HǓ���=7��2AQz?=a��T>>� ֋�?7�|�C�;O;F��nQ�nEfI�T8�-��%1�m�4��hZ��M"s�J<�[۲U��e�xEv|��k�N�m�v�ɲH\�j��X̮���\1Է�<��ֱ�	�[�=Ajw+PlD��Q�I(�B��}-��.��`@tJ����3f�ζg;��I'��sts�NCE"v��l2�s��i1�4u�����{=g��=�i�\���4�N�ʌ&]�m0-���D�`J&������P9,�pc�H,�F�kRhP�Ϛ��XP�����o焺�X�(^��Z@�ֻ�)-�ձ�tC��WgYJՀ�;s��v�p+�%C�ݒGw12�Z(I�_���\��a:v� �N[�����N�Wv�>�qo�&��[kN�3�d��#{n��:{��X'�)�y!R�\�5���P���ИJ���Cn�St�e���@x��j���=L+�|l���~���u��~5t���_�<�z�j*���fD�e$ߟξ��yIr3a��S$B�@:����.O�0v���HO�S�)�H���Gby�v ̽cG��aH�.��G�zƏ�˞����.M�
�z�IU��"OvI�;�C���>5!.AT8��G���2���g$�
Y�g�d���1�W~�۷5K~И[c�G��WCU67z=)�ɐ��A�����}��PVڈ�w0��W��^D�iz.#.��P�튒�-�>G���0L��}$fm ��`}���l[�[�*������}@B� �C"�|%1}Qd���/@=�L�ILr~��Wc�[U�m��V���D�I ����,�J+u��1o=���DX��d
���֙J��t�s���𲹾�N)�����qC�!K?ڴ(hB�����s䔙��.=\s�_�a�`��A�/j����XY��1hq��X�aUMbw���4(aң�C�1���ag�}�i]+n؟P:�@�jf������(6'�R����PC�AJ���� �����Wv)� #�>2��3� P�'X�	�YX�p��;`������OP��Y��v�`�g������C6O�w괰�ĜQ�ɺس�熸���)a�|��rr�l�*�����)Dl�z���=��L�CZ��z����&�
e
oM���pzg�u6;���J]���+�=4�|׷�擅�v�?3�)8^�b���F�qF���c��a5���Va��jPb��H�ݿ*�nf�(�.T0���yr�u�(��>�OŽ��"���>��2Z���\�8������N�t΃�VȑފZ# �g��c;Ԙ��ʀ
�����P�j�_��c�+�&�q�>җ8G�: B�YR�8��,b63�=�}a�>�)�ξ><��:x-A�SV$Z84bT�y|�}��-{#v�
�4Z��W���n�݌�(N���f�_�C����B�OD[	H>�Z���ļ������9�D8��>��3�]��f��,���ނ�fz�j{O��������e�X
�bod:�7���o4pj>��4*��m��fO���]��;�����yBp'ю8�E�]�I���5��lN>�kΚ��3��q����Q1O@w�8�И6$!�A ��E�f�%P��������������Ra�!u�m ���[@�i�E����-���\�uyG\�h�a�S���?]�>
6�|����9&�]�r]��5f�nBCTГ���N)<����t��'�E��Dup�;�FIng5CԚ�����k���w�l�d�"��ɪ�?D�'"�w�2߽g���:�| ��"{#��
�����dEn7q��	t�A̝��ν6�����g���P��q�H�&���.f��B�>���\j/��9���a�z�A��A�X�-��"^�[A�B��W��l9!���yMsu��� �,K��5���<4�6���x+��b�R�ۛ��й��'y�ݍ�p�c/�$�^4��3l�2]��ĂY��+�^���A d
�s2b�Cuaa���	�z%��:Utvx_��d�RvɁ]�&