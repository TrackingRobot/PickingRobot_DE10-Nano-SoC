��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�hF�|��4��פE�5�AY������E-%��T����L*�*�C&б��]��S$�Sv3��X�oq*3���ƀ{y�Wprf�q��ó?����s�wȖ'�m`b�6�eׇ�O�D��#��8I.�'��S���\�9�����_�u�-�9k�^c�K{.� ��Ù�]�"	0��3�=��y}{]�:G`�t	)�GfD�Np����1��?��9'�z�(Zi�Y~M,HWG��p%��be�1b�q(�\KA�C��M���_3%�*sQ.�I�^M��d���-�� ��g���a.<�%�q�4���������ǂ
ܟ���h���:��{F*~ʦ[��G���)�յ-����F5�N�ڔE�F��&�� ��CO=;�d$�r?k����}a.��Pݒ1�ˮ�1j�M*(J�_�IS������gN|��A*���l�-�ۇ!�+��*P^��i";TM��N��BBqkU(���戃rk�u���T4��u��j��`��	91�鸀n�G�J��Gb�d���ź�j�?e�=7�!�W��w-`���J�Z+꧰��s�F�  �%�>[OI|x����HI���%B������mqρ��Xov�#���y��TA�b����M�k�{;@벹�6C&8� f�'�/��>8����Nƨ�ݹ�{��Z�V� �����9%K%(X��$��}=���,߅���c>�E��ge���B����E��US0�|<�6�@ʺm 4'P�E/�Rr)�ŀ�L#�RX�~T	�grI��0s�m��j��O�pa�b<hY_�]0Yķ��;㬭b���vp�m��:\Έ�bj��F�02���-.���Ǖ�|>䦺,��d�3�+0��{��kH��p9�n������ oS+Eu�~Z"Þ0��|NV7q��HD��#c���їщE�g�Yu���%���[sB�@A�*}�y�4��걮r�͏�Ozx��$j�Y����_���3�B|o����,�)��R#��(����?����ȝ�М`�稱����ݓ�`D�PFXh���SU9��~���}m�-:C��c	R$�p�L��$e=R�����'��(���"T[�ף��m�;c^r7fyX���D�H1l-�-�U���Q5���b��p��e�(dxP��7���s�Eڷ���J�FjO�"���R]16�̄(W��eⱱ�$#{�ёu��������� 	���Yy���T��mlV O�Ye��uzb�;�IMކ\U��Q#���r�]��;��Y��@"g��	�����K���x�m탪���Э)�8v[/4��5Rz&����q+|.��u�ۇ ����V����-�d�c96m8�Kt::p�G9�/=!/�k>��ph�PF�=P>)��)~F}7߈7���ʸ(4�+f2��e�*	S40 \�0�X��.���T ˶��v������b5�'���vRf�b���[��k:p����*g|x>�i@��)��a�ٰTX.����u�^��gnr#*T�7��������VP��j�TK5X����W���5����c�����
��1U�n�ޖ���3݆g� �O{?�nv���m�.d�J�_�i�f�~`�%���G�>a0�%P��]b3
�cf��כ�����E�quPhj��=� �m�7��:[֪�`�Pv�����X6א�Ʃ�ܑHO}�o��l�6���ո�'�����(���Իm���Z���Z�J�Q����ec%9�T�����6�x˨�^�!�(�Y��<p�����f��TY�:��q����8+}7��у���yP'ܿ�?ߏF��߼��@�ڋpx��Q@rt�Y��\���#�fW<%��+<���3pM��jZ�0i�]��wY�jn��w�¬qgC�a^`�� -���*_k���jr�̄ 3Y"����)F�[�+v�j��R&0�&���<��Zy�V� �ܑ���f��X�ǩL�L�qS�.��Ѵ<	��1�������+�Fs����*O����g<+h8���v���S�};[�����U8�f+�z�j?��f��a��;Q�4����p�dX���a�e�
7���h�i}ݶ� $׫�R����C9����8����HC&����%��Ϣ��ey��7҆�(y�\ɨ`�6@lY��@<����nk�������G�	c�N�.D��!I[���a2����.�=�E�ɻ�<��&��{��H����Pnrk�j��.L5��Jȧ�gp���:|�j^H���G;��0�sV��:2��o�
}
�r�Y�v�$򴻾���U��5�p|8��EV��'���`��p>��c�>��"-�]����B�7���4\��HACg]��;��EW��@�+d�&����F���U�w�?,���4}H�HZ|\*b������#��1µ�n8������(�o|�G��D�b�q>N���d�O���;Y9+����+�ژN����?Lc	H��m���l9���w^#���*����G���~QY��*4U���O�v�0dM�J�����[���fX�o���v;l�I.��&�S��g��o��������rYX����_��P�݌!8��+���>:]������;���1*R�[j��őpZ -w���N��4�w?8 �D3[��X(ۼ���^�Uا,�d��AO��#u<Y۞�b�������`�)XF��uB0��@A�8L��o3b���S�Պ�-l�����B��6�+NTN&�E+d�&
y~=�Q����tH�;