��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�R_酎�����U`������p�y&J�?ق`gk�=7ටsNG�U �+S�s�� ��\��|.R�����:��)XM��C� *�̩�h�8-���{>��T,J����Gx��j�mv���, ڼy�w���Wt�I^ �{����FحU����@Leg���V=��.b,S��['�#��?zQ�m�%Ly��D`2�체`��z���uZ�۫�Q�-:�%�`��n��B#���x#����]@_��8[4�l��L+��Q��|k��ݢ����i�SHdԸ-�l�����R0moi�ɖ�W@����#��.��?���g�V$�#��`��X54����BY�im�L��{��O�,�
7r���̰~�D�[!����Ԁ��w�2���=��2pN_�?��U��h*"b���E)���#���+;����K�AMbԱ@��ɚ�ø �R���;�hs	`��K�jP�0���׶�=#�����M+���@�\�[�rm'q��=���`t�H9%�S}�73���bz[�]c��9��M�9��p"�s,�S�(\)��Lt�@?zY��r����bN�7S/��QS|�pb��a�ϝ�x2�BQf�Y�]��O�� Ztq��Q�J:J�^�ԉ��ݱLT�hK
R�����>ux@A~���ھٞ}�r��|P8��P_�ɸV_�F,��,�Y��f��]ʦR���W��>�R,�hPwf��{���ko���f��K�H]T��߹MH=\���u�>̱}����Q7�����p�|�f�h�;��*�&�n1��� ڿi���%3۸� �3�h��ԓ��mԪ�bŞ&��ݖ��F;K"�;$�9�g��Ԡs���<,� �}�Κ) ���r�S��b����Ч��Kc\<��^�7���m+7���!�݊�*HW�$�j�ػ%�S��uP�A������G)���k��}W�4U�]�L�q�.n[c�ݭ�'�\�I҇����Ɋ��L�	� �<�@���~͢�Q�������X�����%:�v��Э.L�g�r�c���u\nϿa������l�1���i�y=��fc�s�G��ZA/��J�"]��12�#?�ٝ#k���r��Ȟ���C�nG;F55��mZ�Ջ�ـ��HާYE,Ƌ��H�7��W���箛���Pg��!4�8o�̱a���5N�M�wE�M�j�F��
��2�^�`�o�C#9 N�-e���@��<W�����$���d�-n�=��
%���)+fqվ�w��r��HqM�^��G�n�,�7��U�VRҺ��TX���0�V=d��q��c4A�j��'���}TF��Ƣg�M��9��}�iɍh���YDpp�<S�rt�k�����$�MQ��{.�Y��}��g���[w�%a�aȷ~~�"@,�q�ym�N�sQC  �th	0�G�
X,.pI�R�s��y].�hjN鷗J	�M�=l�*��N����TWJ�M�>W�=�\�cjs�!�%o����5�A��&�����]t��v����z>��Dtٓ��VO2�۬\< `C{��|�(Bxti��XuM��_|�$��%Y�u@{��Z�&J���kzc�Æd��y���	nt���}�qy�~�b���+���G5
������]���/a�ǩ;y���7d�6��d���e]T���<29�r\ށ�+�j*�1%Įq]���RF<�_���+8�>���
;���Ti3��[M���޺�������7z�O�ٍF��z��[3D���in}-φU�L�4ϳ�!�ۆ|U�ݸ���E���\ɫ���+�]m��+M��N����K�k�B�]��g��q��39-�ГX_@!.|��$+�X�~<�mӧv<�g�=<:f�C�|�����I�%}MO��_CxȦw��ߩ���I�M��}%]�'x�[r+�/㓇͒T�X�v xZ�8tg�\b8k�6���l����a\�N�F�� "�-��Y�N*�1Ĝu<���)�rGz���p��6X�^Bt�ނ�D5�뗔��/a��.��XtcNk4S{p���3���E>1��e�1�Γ}�o���8�e+7���g�QO������7Mސv��-�s�����(/���$�����X$�[� ��Ygao%�x�F��y�)x�M&R:��c�z_���i�fˤФ��^�ր�5�j.��/��Q�w.�V��Y>�Os�T
R�#a��8����G�����I��(xev��J�]��'�1����I��s�
����7�]g5��n𨴒��"��vā�\iM"�'D���-�^�M��UBv|�6��2�,V�r��ϿS1]�U���%��������	� �L5B,��Ͽk�}m ͜u��� �+6K:�$�fݓXF���/��
��1h�~��#q\�f����oF�8����$�nFyw\3U���I�sq�͇6�G������[��������q���⸖�xQ|��@�l���Э��Q���^fА��J2���D�h�2P����G������NF��ļ���e�NBd�����Dc�p�m·��3�䄶�9���B�J�Ŕ���jq8>{q���Q��r6���X,��k�:��2S��NׯȘ�. !����t�[6㗘��<�a$�?\�\�b����!���_�'}��[-�{ķf3��S
�q���{��s��#��6l���=�X���Q��i��G�KF�y��+q~��{A�7���ŽH��3����8�h���)���p<�+�G^�%_�:�%x�ոֵb�qkݡ�tᇏ=��+gF�k�E�8�WJ/�y�D�h�L�>Z�{g�"5T��=�]���Ë�'���0So�0	��\�)�ǫw^A�k�ی'ٯ	[�y��ƛϋ���B���!q�&n����ܬIa����r-$o'��VA��a�6��qd��a���C,�qh@�X��P��6W��]$�7CH�x��
�lmC<ݨ��)�t����
���s~��r��lS�`<�N��ҡ��,�!�!���(᝭H��KYAI��� �{�1�$iFG��:J$�*]�wOI=��Jz�0q0$j�;��HW�Ê��|�Uo�O����J��<�{Xw%�ZuF�>��BUX��������0�CF���a!گ`�c��M��,6&0� �!��}m����f��}G����=�&�g-�����v
?�Dد���,m�C��i�:\�I�w�S<�+Ov�؈��1d0)<�|��N�Օீ�D��'y3��s����n�Z3�b ���)$~�x���F|��b�<1��p�dr�ҝ�ur���}����8�c��8颇�͆�Z�:�~{˫�Pū��!/텕H��dx�u�79���\>F��My���"�x���?{���5D��L%�����N�nF%��l�1סT��g6KZr+�^*`�{�33��C���F�����K�GU��Q����x[��^�$�I@t�[������WČ_#��9r��6�v�F*�<�vs�rD`jO�7���r��8���[��W�R�P��2�\Rb��]���U�7�ܩ#:D��Q������چ�x��i�����Ua$ie�<S��8�d����)��k���K$��Q\�`>T�����T]�n�մ^hj�����c�L����%�w�"J�odX���%c��k�7������+�3���:���Iqk=XL����E�0�]��}��i>>/zr�������������C�����4� S: ���x�Z�22�h|��GBL�ʏ�=\5\�������n�=oY�ӻ�O�A�?�Ac�¢V?k���7s�Z��?�X�a��^S]���:w�X��c�`�c��,eCs�^D�� �*2@vv_�F\��Q��RM���G�
8��&#���~�4vEU(�N�do0��mN�)E��bѝh����ڣ�qTLZ�-��<��!��z�+-��v��xA	!�>*�d��km��XJX�"��!o�]� 7��ݍ�	B�+j.�̛M���B�j��� �tq���^����9�Z#L�I����yB������)��k�3_�<dU�A��l��Ľm�4l��)UzN]�x�ˇNU��[�OO�+�&��Y6*������Υܹ���kc����c�$�?��R������)�f����a�H�-\���J���������F�S�E�<���Z(x)"�R`��r���
p��4��ӗ�s��э��<�3��t��o�= [D��ٜ�œ�^r*�x҂e�j�&g�s�I�>��H����&d6� ��џd�FZ�a�������ť<����/%>�oBkx �N͒��O|P��=��#��-^ۇ)�>�����E1 {��f:��m_D��!�-��7>rfѭ���NmN[��C}1��))ΖnqF
�揅�"�.U6���0+��~/�@�������>�'�;w&��<g�#�}U�3��_�f��f�_v�k��䐀�<,6�qOs�F��Dç�/��s�X�R��[vk"\ʍ�Ê*�6Z�7�-�e�vck��9"�}��炥�(7��QI��豨,k~�Ba�lr���-W�`X��:�#�R�oȑ�ɰ�['�*�A��m�M��a�<m{on;��]�:�vbz�-��[\��+Q�SZp����<�8a	����'�}r�}|����u��X��r����Ќ/ku�(
J�&�l�i�R��m2���Mb�����Q��\pYF!6�;�]�/��G��
�;����sL�I9j咸��.e���Kz r�{�f�\�H��G�.W�{ۓ��8lg<2�ˎ^]�?�(l�%�]�]��;'���u�4�j���_.^�R�gS�^�7Rwh�s8��q�{ńJĭSDę,��'�-έ��5��C�j�x��nXh�F�O���u+e2�-��_�D�ȗ�5N��ޡ�K'懪�1��/�6�=e��
9���C&:���$�;	O.�Z7>�Ae���xP���k�FC��mEl_�*��D�Zmy��eGn[F�2-7�.;�0_H�����Uu��2�]�h]������<g�^�%����^"�Boh�O��t����i "R�ny��Z�:�jy8}�t ���4[��u�	1�9�fwU`��
�X;wslr���}�䧥�C���jKV�I�����y��m#U�@oW���z6[b���X�4ᤀ�E]� 9#�o/[Jn����(H'�~Ĩ�<K[Y���q�.7l�z �[�]��vL�:Z�_k�l���,������!�k�.1қ�+f4��������z�y�N�z�WJ0�$�Z�z�E.gb�%��k�݃�2�%������Fګ�Țf�.���(�,&����R����U��);��dt^T�C�8�'(��#F��><I�Eǫx���Q�H���uY��94��5M#�'R�q�����*��[f��R@-ctb�!����L(o*���#+W�BbW�؆�vf"�?�u�@��Q�$(V�F��E�4	bZ��p�ڷ��Wr�F��6��
Z	R�q�(r�,�y�*,���ބ�p�/��-48�:
ƻ����#���$n}F�����[b8x��J�m΢�}��21��l���p~�J$�����}�ق�cɉ�E��	'����!�sGq��6�7�/���u��Uk &�y<
�6���Wz�5��Lm���nN-�����. �_�XF��]�U���]�b�'�-8��a���?߬_D��m0�H&\���p�7�7�
�̘�M��䭈 �|��Y�4�_'���K��Ղ������\*�K�%� �8a�
rF;Go��Q#0��>�Y���gLB�4� �~'���]g��yt�	��+WeR�ئ@�����3�b��;.K�nT�����$�"k
�]�ۮ��~2	_���V- 2���KMy��N������WϞ��7o���;+s���d֘��cf,zxy�uC�)9�k���Xr��>��~�����٤$�i�����LU�[���l^��zeY��N��N�{��7��x���#���f[��<S��9OxJ.0�x�J��I�����N�������J���*g����$}[�]2�?ы\���@22N�"�Hə
>�y��5##��M�*��c0�*���V��)A�h2~m�Գ�cp��z�a�`�9���T#�U�ϝ=`* �l�!��T�����M7MĀp=�*�i�Uu\��H��m�}�����Him�r�#�%}[sw5�����X���:`���~k���y���/d׽�C��Z����?i8EV���M���c��Y�iF�93�l�];�y��Ǌ��ż�W��,�m�N�cӶ�q�De���z��KL�9,���]M� O��J	�ދ���L�H��4�M���޸e�y�/�3��T(�p���|5^��V�ܝ/H��K�cW�GEl��=�	��.��=� ^+Ň��=zj$�j�F�_��Ԛ��/�&l3G�,�����N�~Yt'&�wVH.�;�d�;/� �'��9���C��F1�dF.�~Pє�w��sLw[m	zw$���L�����Kf9��t��r3q��\f�,�ɑ�o��z�~B۫Ut�]
B5���aT%
�+����t���u/x�������q;�����xUH�u�)2�����l���O���o`�U^�Q�ܝ� Pz| �����2)Nɔ`�w���bڗ0�������m�tܔ�F���@F�4uXi��xW_�@��u��8�҂���@'"�<Rn�R&�����eP�}̾��Jk�Z��^�eW��ꬒ�wz+E)��F�HR�1q�ͷ�E������F jZC�h>7�(�M�F3��zUmD���4�����ŭ�Ȇ�^���_R��O^����Dp���suK#!���aqފ ��ك%)�(���ݩ��\-�W���[�LY�Oio���bA*,�_���`��<�Y�2��u��c��'�7�u���?J�D�-�m��	X  ��8s9,���c�J�p.ְ�>��Z�����}a���$�"q"o\˭����ּ �З���
���瀿2���*�X�^y��r����7{����#���������L��S����W-b�v�9����s����2�9㉷��qO��6�](�+��hڶ�����
���F|b�.x =hH7�3?,��ʇ끹W�U\!k��A:�^0Tj�8�J�y4R��Qyd����:g@6�IP�8�*�{ 7҄}��E���'�<.I�>��]�j��a� ܏�i�V#Mv��-��g?)���|E�	���ZsE�c���"���*�G&��{���'&~���(��~W@�

�|eo>Մ���m���D�:�ɾH�M��s���FX�!�ȗ+��ؐ�i~�P�3�K���\xp�3n��ΥE7���8o��)T@��N�	{8XJv��}r6@v�M3hQX�e=sd���1In�T��[I�\vxH�B�}�(N��𑔼&����mkh�M˛�8S��P�vFg�q�i=�u��!�7v^��ŽH'<��Y���s���P�S��d&�_b���ħ_���%;�[͸��'0'�8	�>1���b�q|5�.&���sQ�ǻ��4@ۤ5Pc��������p/�@�ߩ���G?b9��7���%�X�$\���!pe㖞d�Gڟ�F�[+�xj���5B0�M����t�� �?}Fm;)T�|��,�R�����:L��]Iy��h�0��*��qX���ſv�x��)�a���Y@Aڒ����'�v��M�wP�R�	*]9Ay�~��{��g��I����*�D��?�l��j�-2,H=��9��ɡ��=�;�S�d�XLAaڍb ζ'i�<#ԍ"��S��5���. *�l�VL3�;5&!�IM�ݤ�\�Ț���w���/�:Ь�^3䅗�܇W�.ja�d��V�7�������,C���
��Jr�/`�ض9���T]�<�#�>��=��Cس(A��b�c���j	��yȳ�C���W)�zP���ӕŒ\+o9�f��k��:��.�Kl�-��2�v��0 ��#˶�6���N������S0%�*e8�uf6���Mb۶ .�&ٲ��n�Kx������B��(g�0%�Љ����Z
;qin��|n¬<e��K�����@����bW�J���f����i���$�Arհ=*k���lcM�&��H�V';t!ܶ��<�|N�e���UA����B9���c9���<M�٘�%��n���]���v	����7%.5�ިQ�������!	�z��n��Z��(�!��1u�1��� Ӥn��JJ�*TR��l�!>�2�Z�-��I��p "���6��@�۰�%��ǥٌ^�"��c�T
�YO_�pi"DA�J�p� T��ɢ�G�o�VB�T®�5����мX
u���P,a���7Lq������ɵO���zUl���(#�e�,�1,�eB��(^�?���I�����=��^M��dB���-ŇҴvE�p����c����ƶ_�M�����|#�I������a}�!w%s�!���?�ݣ�&h.ʚ�Q��Kz���X��k~J>��D����M�?�_iL��Ma�N��[�;Q�=l6��"��0�3�W�%�W�H<T��''��a$e�{����ć��m{��ȭ6~�C?^y�z���P7�ؿ�p/"�^�o������T��=��E���K"A��[U�ݟ��V�l��'�iX�Y�27\!����a�.{�;�]ȯj���r�����^�����Q�W��8B[��9�Ji����Q��us�D �h����D���$���FܞV��l��dڀC3,�|f��w=�
�����+o��P�8_�0�yr�e��.C͹kT |�iRER=�։ ��Ӆ(@ KnyQ҄
of����6~�u��Z����G�"uZ5B��r�K�&�®'�-*�d��p�_AW����8�$�)~� �p�d=��0T�Ej�.p�2fu���^ё}>��P����������gZ�I����+����C���ԅU��j!��'����|��ec�ʍ���>e�o����Cj;��h������BG��N��|u�5HέQ�?m��^IKb,ѱu�"t~�>���������">F[|NQМ��l�P2���ƏNP��l
�Aw[�v���Fߋ	8D�6?��K����jH���������29	9�P%8wz�+��a�M��N2�V0��	��V]}�<M������-f���*�s�vl��<�D�g/0/�ř+��D]�)��Z� �"�p]�|^��Ӱ]��1[F%s����`��� ̏���t9��cq!q�٭����Oc�(o����ILxY���� �>u���63k��P������2�$H4��ۗ��D��Ûh���]�`M��?8&��5` !?|���a�e�}Y�9�t�W�~�Y���5���x�{����1d�#{�V�.R&�Z�P�RGO���*6>�ȿ��Vu�W�/y����s0�S�s^d���+%�Z���A������~8()8N"�OJg�m@;��,��&������9��|n2-8��,��lHk�����:T������S_�S/6m����@���m�Wg]zބ����M�k3Z��v��un��$��"%R�乼8����{�|�{h��8�jŶ�4�p�^�cVC �}���C�D}&��6�St^a�_i13�<1�١�y��3h��BTE.Ȋ>��3�C
���
���!X����ax:௷�:G�L*��m���6;O)��Lx<c}�5�4�� �gv�%�+-G���2R�;e�2���Q����7xb��t�}
v>�.lSB���b=���Oe�Ѱl"�����1�N2PsB�����$�`��z�O�*�,Nt	_�O͗(�$"8���3��"c�#�6�A�E�{Th`���	lx�EI�W٠�x�P��F���WKG�s!�)Fl���y���+D�����!�f�3T�V� ��1
2�[uw�Eo�/���<��ؚ�����^�_�4�������D*�p�)���x�k�GOM�����c�q��z�O��Ơ=7��)���,�m�z
����r��Q,��f��廆�T�3&�Aql�m��.V'���h�H���y�9�߯�/[�-	Oïa�jH��i]����L�N*�
WMy"����<m�����¦�S]�c[���U� A�2��eR���Z����b�ml�t+�
M��!�;�2���OS�G�մ�&s�`���������{�?������כ)��[q���\j8��y��C�'R��ﲡ��>0�Hay�e/�A�哯�5*'F��f%2�;c��� �S�S�>��	kk��.�W�ͷI�Si�u�`Y�ۇ���~�#;��+���6��c�;�Y(���a����)���]"j����� �c��Sŧ0E���\�WE/y�]G@ó5K&��c1��lwJe�?V����a�/ҝ�%��ث5�^���ۙTJ�8����
3��s[9�`��C��-�3���Y�@c�)�R���Ԛeу�&�qI�U?8��%JD���k�ό��%%�w�8�-�)m�Z��5[��I�S���*�k/���{�`���VXc<-��ͬH)t����s� XhN���ʹ�m�у��������G�Y�W�1�P?{�.Ҹ�E���V��-/#���~�ej�!��� �/Φ!g�H�j�W>�s���ls�%�7�^�k^kҬl����~SKg9n�1�63+�Qc���:�A$A��Զ��4� n'�Y?r[�4��5c��wk'Đ1k4�'R�����	e� �KCfM|P��*D�L�A_Q�{S\�Qp>���2n�0Z��x�D�f�r�	���n,��N�q���-P�b���:���ʓ�s5��bW�s���{m��B
���FV���
�qJ������i�H�.�'F�|CQ��H�>���?�t�Y��규�t
��L0������S�}��U� ȕ2��.`�7P�x��"\��oq�|��@/`z����Zgh�ڙ�Ւ�_���Vd�� q��\��\}�)�qI���G�U�|kA��o �S�����%C����'Y�������5;��zC:�^#Ƙ>5����f%Ǎ�_�����3��[����������س ƥ2�\
����~�LH���^���yZ��~��XH�f�~�D@�.웇���|�Ict���
����k��A3��J�Jt����q&�)ei�}_�)��[� ~|��^�d�B��g�j�=a]�^�MR��[�c�*��s^ff��`A����?���'�G��r7�)R44��i��Z�j��P�E�[?���h%KMsk���٣��ԉ!F��AH=Z>Ƭ4X"ً��j�R�(���ʼ��>�e��NT��ΡD�燛��%�E�����o��.ӻ_�Ҥ�4�-����~�g��)�{@�7y%l�w6�p뙥�h�J����f|�^�F�y��cFN��+�u���ם�~{��
v�<�r����$�p�wE� ֞P%����:''+���Y�6'#�~z4���?DM��/Gϧ�|a_aKӸB�!�@a�D��FXG��V8��:����x�
��YO��­*�]�NpC��B��vƫ�]C���� �*�X���\<���)������>�$���jg&,y ���D^��_����~�yB�8��T[����h���'G��_��J��$������=Ɯ/wC�"�?.9�Z���O54�<�X' ���*�w�C��(N�@�n���{���H2�B����[��y��r���'/�ٜp/��:���cE�a�PB���f�7&Q�
b� |!����k%��F�ϑ��:/�FǶ��[܏����p�z �n`h���̀��\�y�pΒ�MF3�0��"���[3�
jS����F ���+����zU��U����q��0�dh��CZ�D[�܀/������C��٦g�a2 ��uZ�҄����.|�l�z_�(�������Q=��J+���0���1g����������j��6#;><�<a���Cg_��<���}�SN�����YK�������io�3����T��+;#@A�|�&������!�n�7�ܙC_�`ʂ"����G&������`�y�<��D�g�ע{�eh�\ׯ�b������id�%�Y�mX:�,8�����=�eϠ�;���.�C�ʋ8/n�ƅr14DS�Ҷ&��ՙ~A�vV�\�5F�9֌C<�Sp"�?V(���<V��	}n��Y)l��{-�|{���8����t���4k��@�@[�
��3��j���g��_���0MM/��z?-����!�t26��w8Ӽ -	��t\��Vu�Ll�%O-	�yi��
$Y?1�1��|Պ���K�/���U��2(`�yFɛ�/���*���#�_	F���e%3s��S'���e3�	��eßn3gw�FL_k��{����:e����7�8�1����*K���(����)�wҧ_;!ԭ�x�����ꑭ�
�4�l��5fm�5Y;���*�g]������?0�Q�_�4�}p:����jU�\���`�Nr}Vv�*36��y���P:	f��ɖ~v�L�(3'��JC����>�^*�a�6 �]����5���os�<�Q��k3G�2XTB��N�a�7�C�M9Y����g�u�6�9i2���l[x��ߢ�_��!D;L�E( ;�0�O���Z��N*��-�)�C�F�����a?)��[���7	�K�T9����1q�A噷����
����Ut���A�-��1V(ձ38�N7���fo���9L�Ait1V#)��ڜ(B!���<I$p)��s�-�싏��lHx"àZ�f����;��!���Aζ_%/0d�IH��[�4?�B2�x'�ym�b`%g&�dq ;y�$*���=��睼�$�B��!��̙`��ܙ�̰�D�T���(�lQ0��w[���2�K��2Ar=�Onw���i\��>�����'Q(y(�H~��e׈�ی�T��?R�B��վ&�J.ȂD��t8�t��J �į�ӥ��!D���ӣ���q�8��\�y��4i�� �����jU���b�5��M���u��V�]+�/(�U�G�#m�$�qur�t�ȭ�C�m̳�j�B���6�[��!�O��nZ��Bm�^о)
xDy{z���rE��Y<	9r�H��;����n���""���_�@2���:D�]�B�@�(
�t��V^	�6���%5fO�~����]���Sly 6�wT�29�Vv4]'w5^ W��<���q�?�v��Ygh��Āo�~v^n2��S�BD#�ڪ?�ۈ+<v���PZ�dX�'V`�b0���f�+���H� P���\�^�H�\���Y�:wh6�%%9TE	��+W�lH��e�@b��0��SZ&��UGk���y��p<Qi�a6Q��o�M�C��h�ް��O��75g�����ɿ���mK(w	'�L�Ɂ�_�1[p�^'�d�w�C&��D�_t���s%�w�  �y>�	^ʲt����UTϻ�h.��ˏ��W�a�O[�����z݉��Ӄ��cL��-�DU�hhrH5��j��"�k��� ���}T�qj���|Lؘ���Ë �G�請�)�n�r�����5_�V�^�6����|��t=��7�ir�V�X� p�����bw-��޹jˈ����DƣY�ũG���"����2�KN����>��CtL�8]����3��U�Q0�W�.S�g��'���x�
�<�/lw����A���u���Vl���v;��,�k	[�_4v�x/<�B�a�6�ҘH<��I#Ec���3�r��H
e6lW��tA�e�"�3�0�툵���~-�`2�����"�%����y�o�;�6X9�Nz�@�R�K�x���Z�� &�
r������`j�u��s�x-���j�������i�A}7�X�п?2Q�2������~f|������/�;���x��^��gCܵX���Ld��S�� �?F�v��g�[��j����<T���&���Yʫ�~&V+*�>�v�9[b�W퉇Y H�>h%v M<9f��"]�<��K+u.�dd\k�A��v;�E�D��4�_u(	�������W�9$���
���-k���w�&l����)[p9�]�.+�!�4۹�v���/��g�	��窄�*��5xsvj���58�� �+������i�+�9������pԺ7��5BɈ����+� ��?�G��,���S]��|Rf�l�B���F^*ЈK����aq9/~��M��E�@�	:�p������	���#Ǐy<�<O�2w�C�ǧ2௄�C�,q=�9:ހ@�p����,)P��U���yC�����ta�A7�C8��(���y'D�q��m���T�y��
�C�%��J�D8¦0������˂��d-��J�Y��ɚ�5��}꧁��_M.�٩�&l��jG-�z���^R�����CР�F�,s�%�0r㞃2����srKBI%M��}��dS��1k�`ѫB�h8��o�!��MU"�p�pYձ"nK��y��+�f��/��gs�*��ag~{�T�������b���Q
y�8>���W�'�p����A���V��� P��,x��� �\���+�a;ڏ��Ev�ʮ��W X�/19�� f�
�:�{i��(AގFzl"�W?�ٖ�ʲ���9�~�������F�,ub�N�N�y>;�|��73l��i)T��T�k3�RN��~Q
�o�0eـI��L3t|$S�I���+a6^���C>])�l�l�&3?�Ħ�=c6�C^�Pqu�m��a�f#]`S=�G�<B�V1�Ahw�q��wp�qg�T��ː}Aq�N��fp�~Lвk��M�ROɯ{51APfV-��=�nU^�6:q9$�����y"yL�+V�G��~7�@^kp������U��T�@������S��`U��(��dwH�j�WqR&�x����k�� ����o{�1�1)�B4#��8��m]ow�|��y�ꯌ�ܦ){��j`���[f�)W���#�~[qN��*�b���*���q5ɺ�@z��滈�A=�"u��V`�]ڵ�M���O%Ȧ������N �]B�gQv��pb����h��{��&ט�i$��?�\�	��s��utcW�%��^f�'�e�B�JXO�-��l�����x1k���Wd\w�~{��\��]��`VHU���[O7`-nT~kjef�2t���T�	'F�֎x�s3h�>��J���(+�p,���5�q?�c%"�������2�`Y/hA�K���GY�9%���:��`�Md��S�(6��Y�;�&��륮�ejdq%������]݅����g��?�b�u�ȴ�iz%����[k��\�d/��@%/����Cn8<�#8c��b����ec�{�G�|�~�(AA�.[	�>$MҨ][��/���P�L��Is����J�b�L��pO�o�~��J���G� ��y�4w;���KS@O-݊X���80gb)����v���$��+�;U~D��I���"To"o�ֱ�_��3+f�I��<�ǭ��4�cG�\�w@yMQ0DF��,���|̃5��tZ�#%�>\������e�4�iv����+��־R�������v#j�+���.P�@"/ٽ�Nlɩ��A?b�"'�[�u#-�w
w����Ʒ-�T��4�XipU�?�y�m+d^9���˖�_D�؄���7!����6�UhlB������I��z.8�vߗ�����n�g�'�}Z,��V�7ȕ������]�"�7��{�j�g��~o4N��J�*���d� ]�a��*g�Z�<-Y�0d6���B�߷�5�L�å"�!��L��ò,.�{"�E���� ���S��oΨ+��pB#>���[#��j=@�x]����7���r��:c��[WP3�r)�S��t;�
>�~N��w��>�D��з��+����B#����T$4{?��$�\���^�$��\�Gp�a�}�����s���qOs�.�jq�^0���5���ޭ��],U��_�4_����Q���+�p$v��~&9��L�p��J�-�cb�Qp&�Y��Dց���bH�U����ҟR~j���{H�z�(|Ntӗ�ށTp6`+��-q�,Ȩ�(/�=M;Pg�Чp�J��/0�i!^[�d�Տ;.��L�Kh:]Հ����m�͔ݮJVkk�O}c�:�,,�ڢM���+��
e�ɡ ����龻~y�ۘ��{��O&F[������ź����KT��������� ��0Z�2������EHX��ψ|�rZ��*�/ȯ3m(<}L�(�G���ُ�$k�D��,�gNb-`	���FLu�Iӫ�C"�*�?�_�1���܊:Y�)	u�J�24m�r�V����`A��K����4���`BIX̷e���e�H��#`�{�x��x�%&g�74N���Ic}�Ti�Vb������'Qa��Do�������lk��ݽ�K握ہ�U���B�m�s�#��.2��x�#�=�h�ʛe cK�t�$Z4"=��y���.&�{q#� ;	)�m3*!%��ү"�P�k.���a>���Ɵ�&j@>a�/��	|�gY����y��ױ�R*	�+����Y�����o��s�./U�\*�n�PX�l�Q(Qb��P�V]񏹮]����P�~ �őV���b,��&	�;@�_V��&�?-	��Lz©�ظ����7���K��>c�u�'�RaXЃ Xut�`��/����y�kO%6�#��;j�n�"z�bc2���pbj�ֱ���H(}�w�l�� a�'x |���9�����$�α�E�a#��@:�W�vj� cls���L0Jb*9l"U
a�>F��h'���u��p`f���������= �  Sv�cw� v��;�Ε$E	�6!�˨ ?��:5�OT���[L�1�Ug��G��:;j��.=b@�p��56�ޕ�0����d`^��N����?~��.���_� ��,��
I�'�do�)�\h!�j��A�����G={w��M�7�)���<�o��<t8�V� �.����w�*"�J�:�6�<��<,���#�%wk�}���o P�(��E7�XF �qPg��I��Ik;�$,��Sm�ÈӚ�P,�<�����A{L�����V�m�Ij�GL돣s��h� [׀���9}�#��$x�Aک��󐨜4�/8?)��E�Փ����qN�|}{%���4�K2�w<�]^�9߇���oz**�6���])�~�$���kZ�CO���)�tpr�{(���`�,5]�E�u�UT��eI#��![J"q�O��PsߜlJ[��_���Թ���}Uqʲ�t�M�5�[���/���!P�xL��r\�0k�s��N�x��Ł����la���`���Ab�<x)}p����]�:�Mj�%A�ʵfѥ4����a?�Ʈ�@&u{����z��-Ck-�M�˶����9"2�W���-�JI�����K끬o	f�,�� a��4��췓P��?<n��/��=y�<RuW� ���z�@���^F%v�\{���k{Y�]4��
��`�)��]/M��F��G�7u
�W�7�e�q���f�?2NE����ܤ	��糡�[�)�c�࢚�4��_��K��jR)����$��l���.}x��t��\/��@��5ħ��>Gɋ��%�촹��7��q}�i RR�p>�~\��Z�gԴ��t�ů��1@����O=�B�tK4�)���⇃�E�����S�7�Z��E�6-P��EsL��]�:R����j�
�qzê��"����C�ɓ*��Xٰ>�^* ބL��r�j(�Jn�c��]���M�Q;��쭻��k�wxfo1��� W����7ã71Z1���@�u�QΊb��C��QP���9���V�!MA�q�IO(Z!gÐ�������z�~���j����<!F�%��_`QX�e�B���X�dvl����&�5���6�#�d�b��p�-��^"i %P�s���?@��d�z���_��De�B�X�5ü�QNwd��O���y�΅QH	{n>����������y ������Ot��4����\�n�S��c���V�Z!�w+�ؕ�+yΦ�����jQ��0�e�g��z`vM�ԟ5�qn[�_���x��l�ˁ
����/2Y+�{l��b ������pc:W�b�8�����yG��}���4�P�(�HqP���S�mn襁�$$�c��}(dW��-:���7L��������0n6ɾ�����m���^��t+�dUn2{"�;c�QɼL��&Q�!�8۳5�J�����Xɔ�����M��JOP�xS����!	�x�"�����������2w|����F�Ŏ儑��{���)�#��6F��o B��	�C�9��j�	W��¸r�n|��w��賀�`�"��PK���BE�#Ș�l4�}��Z�&~�8�3Y8n��6���]��É��Ê���PX����2�H_���j63d���,��.I�m�����Lݴ���2��
��K�4�>9����A)7D;:8�R1B�m�U�S�H[̦����.�M��I�����ȨO~��K]������,���C��@���jBI��m|��nc�x'΂��]�`��SK1����a��V�U�v*�=� JgCZ�R��jm��E���xb���b��Vp�ȯ�3vN4�IJߠ��EC%&?/�ϩ�)�/�ʂ�G�}~�~���jv�ޗ#8.�Vfi��)B쬇�"���dҮ�5�����nu��@m��	��p0��5����|z[�yb���0�O��%�C5ai�K���bR�m�#lZR�v�P����r�oQ&��v����&�/��J�ʮ<	(�K����6, ּ�o��!�J��7�s�G��D��H���Ř��D�~Hۖ��>Y*�ou5
�!Z��l`�/6ό<� �x\�A�rCM�0�Kg�g�n�2�h����`��E���V���J�i��h�l5Xx��|/M��8G��Mk^+�S��̅IMr؉�I���o֡}��_��]o��8���^��!-�Iaj���M��n����ԕr�ª���0+m)�:���@�~E*V��ג��Z�'�c����T7����Y%P��V5����x���5ׯta;yJ,�AD��6���F^ǲ���L��H3N�O��Ul+���$�=TM%��
�ѯ���c �$>���5c��z���s�\r��zF9 :: Y�2��������v��G
 ΣPi;B��D���'���+���~�x�O�o����=��Ь�����jV{JB&��1f���L:>�h{��CK&�)_ϸ���}J���EW��}��g-f2�//dM���ə�#���w�/�v��X�:>��>֜�7$�$S��_��^�$����Lz�hv�k?�7݆�,G��FO�����S����ۥ�Fj���Hg�7�c�@�<�'L2�J��Zd3axH�L��m�3�-�]��@��MT]�:S�u7�������
5�?��iG�4aOֱ���L�ʀAH8����KX�g�(*����oR���;
�!���
��
�z�N�51�U�Z&1ֆ�n��F�%A�oD)��˺�2�[뻓)�P:A�]���ugp��>����pնT��U��N]�&���-!CcIe>�d���Ɍ�:�9*ˀ��秥]��2V���� h�f8�X���r������rЛ���"C��Iz�/x����n썭����~6��4l>:y����'.0��ܿ'�qt��Z.ɝ�Lw��W1�E�索%IO-d=����?�f��s��az崱����>J�`u8�ڷ%1U`W;9�����\�`P�\Ƒ[,��#rtY
?���,�9��O��^Vx�e<9�Ζn;���V�[�Үj	��GY8?4�ZO�Ґc̥n+d���S^zIXΔ����ӧ�LP���$YP�g������խk%��aqɥ�ǹ��ڮ�+�p|ۯ��%ѼY����\��8���3��~�d�}�Xg�]��O�f�{��A���kȜ��)�hB:t��?���5�WQ��ͨt�*�A�Ө�~��$���霟D��<��IM����X�'7ŀm��[[X�µ& 	8��,V:�^���B�B�d��܎���/��ظ69S3Z��\�[��od7��-K��UB�������jJ��E]	���v}��'��T��mi��k�J��k�]C�0�I�RD��R:	nEz��S�,gI�r&7��1<2]�AK�n�t{��$;�z������)P�c+�@�zǧ�$>5�@�ou�eP�UXU�M��"-`#�r�R)�ј{���t���P��Ay6�3�6��R[�o�uԔ�TGDP���ы3��1w�-g����zZl�S�)�{5-`ד:Ò�J�J~�P���&�@g$�Cr��%������䑂eǌ@��WM�2�xB�����*�'ݑ�ܤr����s�`�L��M"<^��d�q#y
u=jSX
m}uɉ���w���$�$\�Xʂ*�� ^��U���*���X	�^�*O�~J�h('�:Cm|V��j��=��9V����]��NSTn�z�W׭�P�@��U�ڽ5�M�)D�&T�th����C�,��6��(:��4��W��br�2��Z8�(��&���&vW�[^1�jJ�TlKT��'߬��v�]�r��בJUR�	��&}oф���yNz��)��w���FM�N��!
*��Ј,��6b��3�)~���u�J�s��d��J7%�u �CJ�up/��TXhp�ؿ����hm��U`�?���(���Z��k�i���f6�p�.1V`�˸���ybɒׁsW\+=�=l*��ګ.�ǋ|y�;p'Y;��
��
�;������1��"s_��M|N��s��RT)Z�o�����GA��C��?�B�o��������&2f�.���dF�V�җ���������������A>�UR�/#!m�G̸c���z���^�Ԋ���aL����S�z���<)�\:{)���UGg6a�V�z�Î���h���{�D��O��$���Y����~]�D䣡+�	ȞJ��^�M���Kk��E�/W,ޤ����Hݼ*�wt�P|��3�S	��g�A��.����7�_,Q@؃���q����q�!xFd�`����L��h�5����4�D������:�� ��W���bZ��U�0���3�;��!ͥ�YJ(��*2J��o��2�][�����&��FeU����<Uj�9�ɳ �#۵	7�n_�uF�b�h��(�@M$�b���Kބ���=����Acv�"�BE�(�u��ɺʐh���m��2*����Z�<�QZi�-9SK«��e�)̏�2?�&c҄�kU[���&l@X��b<^��d�`U��^��-�H� /M���݇��2��6�pjˢ�()8��Q�SMδf_C��b���Cj��DjHXwm�Z��z�Ch������8��ʛ���������b��دs���q�����x������18>�
I-KE��_J���֜"�q��<����� �A�(��)��4�{"ڈk�&����XƉ��ކ.��l��yY�+ �7B�0yIγ�,��-7y���PSHF�/�:��V�4��+���� ��S�V�¯r"x���.jm�~��I�C����6"��J���:n*��ɕ=b�Ph?���4�T�o�����=�Oi_-C��eB�UZS^�h��8�w������29)G�Wbm�^��<O�j�,`	/&o��{�P�fsQ.nI�	��y�m�?C��2�8�Z��������H��j���H'��H����;Ix��xEя�Us���`�Jε���4V��R1)ȡ6��*�{j��z�
�!7�rU�{"�и}C���5��"��`�a��������A]�:���3
����w*�2�`�U�<tE�C�/��ns�ry$?˷�����e*,}$�lt4��w8��5�I�9(z�&VC"`��?��'6
�C����F�Rm���3��1ت����uc"�������Ij��qoI�P�l��W�Oq�|]l�Q�N�`&��8��r���ٍ��m��늧���w��j� �#�>庍}�ijg�Rt(��6�{��-���G�<f�PQ���
`Kg�w��G`$7���dv�&uH��K�9�@Z�j~�Xb%�l�ɇCe1�N������(Y��Z�	=ĒD�R��4��G�K�����?��B+
K�ٍV<y�N������6r�F�z�c����1|��
q�mw��T�|��t�]f���L�~�<N��y�`�|�M�=��N��ز������/�2z��x.g���Fv�+UڙSb/@�0�d�_�.,���R��|����Xi��s�jA[��?�@Q_�pŠ$.E�m�E<e�A��xJJ����HޠЏ��a�zY܈����f���8ʜBd2���`�ۍnN\b�v*��(Ek���0k�W�=#*@���b>�����P��TZW4�O;E�3���I;hFzk�0JI�c�5f#\פPyJ���UE� OG^��6J�����}��C�QޱDK�+����я0���yV�g������Q�y�ʯ���6 �9n���7���f����S'S�$?UT��R3vUR(ԍ���G��>er>D�-\g���|T7&ɠ�y��]A	 ��T�]
��<�4���)�>!�FԄ����&#�x������Y���$�C~x�1���;��Ɖt��&�->�B��tA�"O
o����O1ѷ��y��&B�����W�O��1ξ��hJ����b����y.F�L��ֺ��-��]�"�:x57v�d�K��I{���;�.H