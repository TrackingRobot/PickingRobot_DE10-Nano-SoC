��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�K�7�jQѣb��6���>!w���a%�R�sßb������?��@�?�����J�F�	�����!��#����q����Q�&[(m�2�,�4_%8�/EQn �����	�~K���94E8�z��#�먖v�rkR��1�[v��N���e��ghk������K�D �[֊���md4���k��v[�r�V��u�q�~FW�%����A�9񸐬�6�$(H�``�3��M,�{ ��-ǒu���������K%���ο��:f<A��,��4�8Y�� +
���@��N����vj[�e�Y���q�z�rBl��M���h��A�1E�I�)&��p�_��(�;���ؕ�e�u̬v����P����.�6�ޞ3�8_ަ.��� `<�����[�}�X����Md�3؇%@����р8 ��#.ʊ�)D �^I���)J��-���
8�E%�C�}�<tB�O�ƥP7�Jk�g��S-w�7y |[`Ņ���>�4��2��Ʊ:]�s�-���G�>��Ƭ��q[���[���;�CY-�M��hn&ǥ��� �N(�q~��0��T�myS5�6�)+Ai�h��2{��y0�tˁ%����-� x��"A��=~�߁��)�D�n��� �apo1Aλ�S� �e�_�)�@w��W	�	W��������I�%#CI�*�O����`�3��]���m��q��~�w�4%Hƈ^�rAT���\����F���ԁ慲Ʊ�&�7�ٓs��
�C� �b(��H��NH��@O��1f�m�Q8�>v�V���Bl�ߑ�����I��zIf7Q� A���"dl�>m�����ܪx�W����(��s��Y����f��m`���֚���ٲ�x��M`����AA����57M`$��3�4M��g��!��Fy����sO�d|�27�J��N�j�a]'A��x��&b8��4�`z{L׎��W�<�2���(�����D��3�Cbv�B�9d���_Չ�p�w8���9��,���.�q:hZ�dv�Ew�ݐ��J,��,`��MW�w��B�f&bQM��'����ܛ��M���W�r4.Á�@w�|Yח*��PE�R���z�m-���� �����tr{B-�(L�0O3����r��?�%u��.D�|�T닲!Y�:�Kx�>�!����{�0�?S���ƒ��ǁ��g���e���ۤ���N�m���^<뻠���/8�.Ju�q�Qz���TF\�l��!��	h*��u��Q�K�P_���d[:��2�'�,�cĩ� :͛����2�l8�Ys:m�헌@�g� u�,� ���f�$j1�i�f�ec��l;�ҿ�Gr��0��?R��	��x���^�_�r��,��,�8����ۡ�'�2�-.�ⱨ(���EzHfx�,*ܶ�����ԟռ��� ��\����Y�B��Tº��+�X߰Y���H�K14W��gV��_ק0��pG��'�N(%�-��!E9���������k��y~�"g�:���E���\�m��5��$��A���v߅�p�ֳd�5|�ӫ�����+��#]*E�Ck�񟵥�?J��=∗�a�574���46e*q�
�g�ZC	'�--�3�x�!6�^hq=��:�R�6΢�>�u�ǦS˃v�8~�en>�KP	�]��4�E�9AZ���S�2� a�����c��^`"���0���f�O�#�]��	Ar[�����j�����3�#/ �97�B7|�R�QVU	x����=����2ʬD�z��b,�t,�ڸ��糋l͕��X�]ᦍ����U����|O���1� Q~BZcb��@��2"
���������ʗ����
� �����/�>�S>K.�� �l�;�/j' ��Ob���M2EZ��wFEX�$�	=yb���L������ߌH2AB��D��í6���d���Ć���2���l�*M|�97�w�.�蠒���j��p�K�!(�s�� ]���鼭=%[}�D/��E���X���]ZQH"��iB��L�	q����fP	�+2��麉�i�V4�_{뷁������;ۨ$��:P���y����-������'��-�Rlc�<�{޾��5nà�ڻq=��I�l��hEǊ�\D�9S��?-.���/a���sZ9'[�?�a�GM@o_���Z�m$�o�k�����F�mwV�� ���V��(l+
�=7`�&�d3�P?�����u�Csdg�	��`80��;���Y�RV�>��0lCZ�%[A�1S����r��{'�We�/�|�@._ކ�7�X<���ҙ 1�;$|U�R&c���^z~�8�tA���ޣ�}�r@m�Ser����FNy�Q ���b�ľ� ~��F�E�GYz-eG\�s��-~�wE�3F��$���[�TО�ڝ��帀tp�h\���̘y�I�eוc�-7�N�� ����#�0�ޠ3���C>|%�v��܈"���#:<��1k�+��Ҡ.�׌��Wf����+�[�g�X*�({��1k8$��I��sL���ѣJ�hG �د�~1��;�E���\8	���<,�,�}�����j�_��r�P(OUڼq��W�a���w-�u�m��{��^\{�<(�>e��;�.��v:��L������ҕ3V�1t�͏$�(����$qP�0O[))��)`i���#���:����9g�; �6�f�cE=`��VG�ֶ\8����
ڍ7���k�h�.���)���u�+��c��k�ZL�.`�5~v.pp�L��4a�2���UL�B<kyg�Fũ i���Y]6���, �����WO�������O�Jቤ�d8���mH��,+��E`��3���.�J��V�����V#ܕ�:^:9i��_�w�*kA��yC|<s���mH�!�����*��T� -�V�L�nAp](D���c���nI���8��[u�5�څ�/0��q��ש�J��b�5�;y��B̰Z�����:.����7�9]_��w���W?�EO��Cݩ9�bg�-�� ���@��� ��+�p��鮮I�,:�HR�K���_r���n�J��A�Ez��]*�~9����6��[��@�a�ԩ<2�4~n�e8�[�d]�l��;�V��@�Aid��uH��g����ɕ���{�:�N�5�u���h$����	��UΤ	���$�8��Q���
.?�����-�a=&�������¤��>��PhH�����6|�7v8f���:)b��A��H�(:<4�Z��,��}�!�@Y*�	H��'�Sz�U;g=�����Zgq�QkC�Wb����a���>�i�Ԗ��z��59Q*�ůQ0Pb��4���@�G��'ޠ�֑J���{7����x�i�٥��=uK��3���Ɨ��\ߗf+`���
�d��I�C���O�������%���u�����&=��@��ڙ��WF.���Pn�d�[���Z8}���}�����`���!j5�p+^�V�T�ǩ��4=��D��3����z��-o����i^�H���5�J�p��@�)-��h��^�?�藰���i���۞������4d1�!ͦ	��d�� �W��<U�pꃲ]*&_͔>>r% �Ȁm(���b��\�J��g�MJS�`�3d�_�ů#��p�Y)R���αAk����1���a9[�8��B<���MQiV�s�~"�|�ý[�<<�8YJ��wv�&5��cm�X�V�l]�X}��1��Ľx>K$7Ρ���?�tSG��Pv�����u�g�Ȫ�1��{��d� %���k�ˉs���~s@��T�m�Q&I�r�s~��q�bCOI	�ܝF�4�%p�	L ��	���Fr`��tt{��6�NCK^��cO�ɊM��]Ŋ|\�miApU�^a����o4&6]L�D��� ���2n1NL�>z��j�IK�=1V���-P1�#�����/�ق4E�(��0�%�t��81j�P���К3�ot7�_�Bp%���RB��m�.����p�(��7%�L�P�06Y*�ix>���>���*ވvdkJ�q�[ο��V1���/�j�P��G�Tݬ:<��x�,��P�4��\��cO�9B�T�9����b������j3�@s9����/ˉ&r[�bW�@�"H`7��Y"�­�F����a��]�a�Ap�p�R��H�5X��&�����3�򛎍�#k�9o<K�O<pME�N[��C��f4�D�f-��	�8�RH�&k����=ck2!�^J����t炡-.�D8���Vűx7n���	���	|@�x�m�X&Z�Hk�:�(FӁ����g�|P��_}g�*�X~S���W�Dɗ^�@��w�l��L��'�D���RX�&���L,�B��ߛ���y��8��)n�5w1jئ�B֘o|x�;s��4��>�]�c�w3(ɞ�^��}���ʤU��VJ)s�����+}��]�i�GX#�(4:箪�JH	�褌΋`��ܗ�\O%��Th&LەmX��P�2�<8%e�3���B�!����c�����f`���m�[F�O�z��:<@�� b��h�T��P;�%d��y�ԋ����n0��K>P��_��-�����J��Ec��J��@��A5�P��1Д�9^Iŕ<9c�-K�f�T���'3=�᮳L�'��&3oP�����;M$����C �F�9�A ��F��c�讵�:�k�ҝ�<
��4��L��A��T�.��nBm��]{G��+�.���n��NG<�<����2Nq>�����[�2= �p���z��V�sFX�sL7�)�a��+�QX"�Qr�Q�>YNϼ�hG1��=(�Ln�c �o�ζurhanzKͤ��D;yV%��͝j��Ĥ��4�H�w6�d+�p|��Q�ԇ��R�Ju��kk��`a輲^`�L{ �-��D��V<�[L��ϓ���DD�	'b��If'�)<�q��c ��P�B�WV�o�r��e{��G����?�G��*�?�Z�%'�G6��[�Ԏ}�GkA�C7���²�ĝm)�y#_t�����ac��6a]�n>�-Lh]��=�Z�{�h3�Qr'VPr�D��z�%05b�O\�g�B�`�M��2�@��JN����4H�<z��z����A[Ϫ'�j�y�Q�F.9l@��,��6P¯�v��-r���G	�?j�H�j���3B�I^"}�����%�z	 (��-N!�*2�ڹ�9riM�������lӨ�g����� 1��Q��}�ݣ�=,�������1d��nLb�����1s��N���~�H�^J��f��g�ƬJ��m�I�����hD��fV��lB�O梍�)�j�����-��@K6j��6Kz�]�E�݉d����H<$��n)�e��
'W�"��Q��k�{TsE\�=�Q��?���9�D`�5���: �_�S��`�ʊA譏vX\<~����h��h�i>���u/�b9��>i�Y�rd5E�M���`'.�^�_�U�5,!:���;�F���4ٝ�S�0�R'lHCi{� kT�A<�������$�Ȭ�R�|D��$
JB,�܃p�?aW)�o���n��B��*-bj�}���0���ƫ��ᇱ9E�?+ �������%ZQ�sN�]B���Oɨ�a�@}ac�O���7����?o���Δ�hGV��6����+`��|������4��Xg���q�<���N^��m�#��O�|Iΰ�?Ö)g=8z���:��Y���&�0�#�e����H�xg�S]5��4�K%�U��LZ�|�|Nn�h����Q+���S(3�3����=�>E��$3O�����ǌ"T_���b'�/� ����#\��w�|C��Bbmɱ�}�!�P�6���� ) V��\�-���~&�rJ~(����@����5`8��9I֩ݫ��-xb��B�%v�q�Gx�mJ��}��Ǿ0JmзMw���w��{���Z٨;N��S�x+B���-B���|����~�k�u�zٴ����<�@/+k6.GE���,pTI�fJ$�Y�}���]v�#�_7N�Fk��j�����3���V4��l_.i5�-�0�袟��n�Uc4��?#Nl�fD�JB����_r
�z~�⚩����XC��ku�I�3S�wz�(E.,׈2�D�
��
�&9H�ً��u��,��۸��W&=]pJ$�#r˞4�<��(�S�#��~����^p���%h�[�Tg��e�VǬ���~dH���-=f0�~ۈ��rY�'��"r���as�!�����i��x8GLG&-��
T���PWD�$��<k��wT'���>�����5c���ֆ�*s9~���	NQו���K�S�|�!�;(]��s��i�$ZD�Vh6D�P���l��^�t+��Q��>����B�Q���۟�ڈ4�HQ<�%�1>������>��^sM��.�kH��NB`7!�_��	�}�����_���>L���*� ����x)�Fmεu)]�������s�F���~��L,`n�hvcF�%�O�Ԋ��lZ�����s�l�ru_-�3d`�Z�y*�ke�O ��{k|��q9�"RU�1�!�!�|��6mEO��u@�x�M���<\o��r���Oe��8eI��`���TƯ�
����H��M�?�WK��sNN���QZ��S@��2C[�9��;t�ѣ������JxW��:ډ�� �(�s���9�Z6��g�w)X�ޠIiP�"��d�k��+�1�n�}HC>e_��m^0qN��f��O����n/��f�"CM����5,�������󴁇k��p ��e)S��"���;�:��oYt��ЗjJ�.�A؁���o<���%iF��K,>�j��%g \y���f��8���\ٱ�w���a@p ��9���|�sYi��k� ��m4f`��]�	+��ue�> $�#�;���-%��y=΍Ł��!X��+�mb�H���'M�I��2)�$�?�9��AM[!Y���Bh̴�N��G������2����Jw���nC�wݩ DTO�Ҩ���`����y�W�[�$�/��M{�_^ދ]��۾�g��h�,U��y@�q@uxu&h�ώ@�1d�5�Q������u��f���Pm�BaT��hG�w|M�D�]aJ[f�p�-�`!a�j�{F�N�v~)�p������_}����N��?�f�(����9'qڀ�_���A#���e��5:�AVK.)'Z&��5����te���H� �V3��!�w��caBs	���o�z����Tڢ��ϒcws�ju��) �{L��;;�d�|.BHk��1�=��� ���e�pa�w6y7�ح�𘻬\���n�%ڡ������pw\x ծm�Ձ�5pA��=W�e�s!n&&���Þ;<s��Z���O��E����W2�$h$���Rf5��r"����7%����'	 �o���a�Ʋnorrt�_���'�ͭ/y�ǽ��/����]�U���F�-��3�[��
�wj��� �*��ŕ3a�y(��{Hj�ĜV�_?���4k���Ρz{�G��
Z|�̕A�w0yXO�XSĎ�����9�yk��Q�/UK��	��I��Uk�bϗ�5�6�w�����T�
���ܥ���s���Bp���.�e�)I�=���������p�_G��1�^S��WH�Q�Ve5�����GCn�M�u�|X��U�8&ȁ�K(s!a{�n�)y�l�����֓��K��y�X�PU���I�>��}�ߙs��$ՒY�P�9��=e�<A��wa:cKX�2s�*�Y�X�����BW)Rc2���s���ì1^K���ֲ�4�xYx"-?��S~��k���r?ٞ����\2l�=~�Q�٫8�f�0�K��{�<���Ѝ���!���/з���ei�@~�d�f"��b�5��G]e�n~&�0��V��_k�&/?����E ��)�Rk;����1@vy�Ƹ�*�NS=�����8�>�s̗g��4-oC�.�����W�S�7�l��gs9l�+���ԔX���D��'�3{��܍�ں�u��,o"��ɸr1�A�5�������{��ڶ뜓��[�L��|��R�m;�w��*欑'�e.�ze<��L�\����(��}E�J}��?�͓k��Rb|��zmo���f�y��:0D�̎&���u�����8�b:t��a!����ʀ9|8�~�� ���҅�Y<ݾ�ix�u$`%��Z;o���Χ�Y��iQ�
A�O�6��"T2���>$����?ud	$��j���ln-;!�UޟGA�Xd���5�-p�ׂ���{9H'�m�}���A�c�@�zvj�'�H����"
n�mez)�^	��
Jo����s�]�o����._-���\n������\�h0 �:)y���?Dhsc� �X,��G���/d�!�T�3���/ÊM����!#8٘T#'��F��g�Ka�($��w���)�H��*@nj� ����A1�c����2S�X�x#b���?�u��c}
��r�H�3-�K%�b���E�
�����\N�e\���c)��$�G�%$��%����^}��i���h�p�ߖGvo��˙^~f��E8@=���R1��Naڪ��]����U�9���{��8�� -�:�:���מ�olA�z5�����9�$$:
�Έ��L ���8�Н�{Tg��X�"+��wv�����Y��r��-��˭�ޞ�g�K�7+���鎕oɬZ���	�o1NJ%5���:h!�N�uP���P�T�/ە�i;i[E���Lz��bz�p 򼬏��*��d��0��vtV�2^l��t
5���:�*�;v��g]t�&��6Ѐ{�����Ur��l�LY�X�(܀�i�A��R$�57AYH]��BL"��e@+	�*�<`��>~����Jӥ#5���\���<���ogTsАm�Є,?L����l���l�Q��n�}��K��rU���m:��fTs��ꄯQWIZ}�&�t�l Y%��PT!�>�;�ƨ;��y�d
�� ~v��{cu�{����a�Ӄ�#����nȂ�.�$\w���m<ak_`�Fe�i3EQ��C�.�/<<���4���9��.Rܙ�����yǦ�U�\��m48�u��%'�*��}�C+>�dB�9������
��,���UK~o������G����=p��C�a�m`y����*�RO'p&��̢�׵���Af�1|2���Ҿ3�u�G��%�ױ�@5�É�捅�����j�|{(�x�'c����q�Iy����vU��q��`��9oF!	���]�?i�����*&�߾���h9��yR%|�@��"X�I��Ղ�������E큢ƯVҤO��u5�ޣI�{\O���d<jo��A}L������8ͥ����l�L�)�J;2-� Ii���*)
�Jod���BB/�O�����]3��NA2�$5���׊������.{~<�w�}Y!��)��z��'������HM��-6��0���[�fL���`�b�ۻ�}�ߡD��g<
�1�wv���� �E�	S>�l�^N���&�:�x�J����Y���Jy>���J�ww�i�Kw�l���C�A������F��_��|d�����Qۑ��b+}�a�kV񿤪��#��mk'�mBב�Gx����N"	Mb�ˍ�<} 0�0]c�n�Ү��cUy5�*��^�ޗt�\�W8���);���_&Ь�WW�mog�=�}�����e\�o����mO�'�FD2�[��ρǓ�P��@Hl#^�H�C����ALpb����G'��;͐u���[YJ���޷H���`H�`����&�s�`�n��:@u��W� vz׎Gy-��壉(�`��.mr���=�u�(�T�/KhX�*��Y����sk�y��G6E5�Q����>����s2['�]K@�40VL;��3�SE�5�w5��D�0�1L~Ɗ�=��M���|"bl���lXVƨ�r�Yt ��t�~O��z'�_�G����[